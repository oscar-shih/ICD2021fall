`timescale 1ns/1ps
`define SIZE 10000
module tb_mode();
	
	wire [3:0] i0, i1, i2, i3, i4;
	wire [3:0] mode;

	reg  [3:0] i0mem[0:`SIZE-1];
	reg  [3:0] i1mem[0:`SIZE-1];
	reg  [3:0] i2mem[0:`SIZE-1];
	reg  [3:0] i3mem[0:`SIZE-1];
	reg  [3:0] i4mem[0:`SIZE-1];
	
	reg  [3:0] modemem[0:`SIZE-1];
	wire  [3:0] ans;
	

	integer i,j,error,error_total,error_part,hide;
	integer err3,err4, err5,err6, err7,err10,err20;
	real time_avg,time_step_sum,time_step,acc,total;

	

	
	mode_max top(						.mode(mode),
										.i0(i0), 
										.i1(i1),
										.i2(i2),
										.i3(i3),
										.i4(i4)
										);
	
	
	initial	begin
		$readmemh("i0.dat", i0mem);
		$readmemh("i1.dat", i1mem);
		$readmemh("i2.dat", i2mem);
		$readmemh("i3.dat", i3mem);
		$readmemh("i4.dat", i4mem);
		$readmemh("golden.dat",modemem);

		
	end
	initial begin
		$fsdbDumpfile("max_mode.fsdb");
		$fsdbDumpvars;
		$fsdbDumpMDA;
	end
	
	initial
	begin
		i = 0;
		err3 = 0;
		err4 = 0;
		err5 = 0;
		err6 = 0;
		err7 = 0;
		err10 = 0;
		err20 = 0;
	end

	assign i0  = i0mem[i];
	assign i1  = i1mem[i];
	assign i2  = i2mem[i];
	assign i3  = i3mem[i];
	assign i4  = i4mem[i];
	
	assign ans = modemem[i];

	always begin
	    #3
		if(ans!==mode)
			err3 = err3 + 1;
		#1
		if(ans!==mode)
			err4 = err4 + 1;
		#1
		if(ans!==mode)
			err5 = err5 + 1;
		#1
		if(ans!==mode)
			err6 = err6 + 1;
		#1
		if(ans!==mode)
			err7 = err7 + 1;
		#1
		if(ans!==mode)
			err10 = err10 + 1;
		#12
		if(ans!==mode)
			err20 = err20 + 1;
		#1
		i = i + 1;
	end
	
	always @(i) begin
		if(i == 10000) begin
		    if(err3 == 0) begin
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;231m░\033[38;5;51;48;5;230m░\033[38;5;109;48;5;247m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;172;48;5;94m░\033[38;5;172;48;5;137m▒\033[38;5;214;48;5;143m▓\033[38;5;80;48;5;254m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;29;48;5;101m▓\033[38;5;208;48;5;173m▒\033[38;5;50;48;5;223m░\033[38;5;138;48;5;239m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▒\033[38;5;129;48;5;137m▒\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;166;48;5;180m░\033[38;5;42;48;5;244m▓\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;86;48;5;101m▓\033[38;5;69;48;5;143m▒\033[38;5;179;48;5;136m▒\033[38;5;130;48;5;173m▒\033[38;5;50;48;5;223m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▒\033[38;5;80;48;5;101m░\033[38;5;94;48;5;95m▒\033[38;5;130;48;5;52m \033[38;5;180;48;5;94m▒\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;94m░\033[38;5;172;48;5;130m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;43;48;5;223m░\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;230m░\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;100m▒\033[38;5;172;48;5;94m▒\033[38;5;215;48;5;52m \033[38;5;172;48;5;94m░\033[38;5;179;48;5;173m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;215m░\033[38;5;172;48;5;216m░\033[38;5;179;48;5;186m░\033[38;5;172;48;5;180m▒\033[38;5;50;48;5;224m░\033[38;5;209;48;5;239m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;238m▓\033[38;5;214;48;5;137m▒\033[38;5;172;48;5;94m░\033[38;5;172;48;5;136m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;216m░\033[38;5;214;48;5;186m░\033[38;5;136;48;5;185m░\033[38;5;136;48;5;185m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;223m░\033[38;5;50;48;5;224m░\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;239m▓\033[38;5;69;48;5;180m░\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;137m▒\033[38;5;172;48;5;58m░\033[38;5;216;48;5;234m \033[38;5;173;48;5;95m▓\033[38;5;208;48;5;137m▓\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;202;48;5;236m▒\033[38;5;208;48;5;95m▓\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;229m \033[38;5;221;48;5;187m▒\033[38;5;87;48;5;230m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;235m▒\033[38;5;50;48;5;187m░\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;186m░\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;95m▒\033[38;5;221;48;5;95m▒\033[38;5;179;48;5;95m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;221m░\033[38;5;94;48;5;221m░\033[38;5;221;48;5;186m░\033[38;5;178;48;5;185m▒\033[38;5;220;48;5;179m▒\033[38;5;220;48;5;186m▒\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;51;48;5;230m░\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;203;48;5;186m░\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;222m░\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;137m▓\033[38;5;179;48;5;95m▒\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;144m▓\033[38;5;221;48;5;230m░\033[38;5;94;48;5;224m░\033[38;5;82;48;5;230m░\033[38;5;131;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;50;48;5;180m░\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;172;48;5;101m▓\033[38;5;209;48;5;232m \033[38;5;52;48;5;16m \033[38;5;209;48;5;232m░\033[38;5;208;48;5;237m▓\033[38;5;136;48;5;187m▒\033[38;5;220;48;5;223m▒\033[38;5;29;48;5;224m░\033[38;5;131;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;220;48;5;180m░\033[38;5;178;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;143m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;144m▓\033[38;5;172;48;5;144m▓\033[38;5;172;48;5;101m▓\033[38;5;172;48;5;238m▓\033[38;5;208;48;5;235m▓\033[38;5;166;48;5;235m▓\033[38;5;172;48;5;239m▓\033[38;5;136;48;5;144m▓\033[38;5;220;48;5;187m▒\033[38;5;42;48;5;223m▒\033[38;5;174;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;207;48;5;180m░\033[38;5;178;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;137m▓\033[38;5;179;48;5;95m▒\033[38;5;179;48;5;58m▒\033[38;5;94;48;5;236m░\033[38;5;136;48;5;235m░\033[38;5;220;48;5;235m░\033[38;5;220;48;5;235m░\033[38;5;220;48;5;238m▒\033[38;5;136;48;5;144m▓\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;223m▒\033[38;5;87;48;5;230m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;88;48;5;232m░\033[38;5;50;48;5;187m░\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;223m░\033[38;5;99;48;5;230m▒\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;80;48;5;187m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;51;48;5;230m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;80;48;5;186m░\033[38;5;220;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;94;48;5;223m░\033[38;5;131;48;5;237m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;50;48;5;186m░\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;222m░\033[38;5;214;48;5;223m░\033[38;5;94;48;5;223m░\033[38;5;87;48;5;224m░\033[38;5;88;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;173;48;5;241m▓\033[38;5;221;48;5;239m▓\033[38;5;43;48;5;180m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;178;48;5;179m▒\033[38;5;220;48;5;179m▒\033[38;5;69;48;5;180m░\033[38;5;50;48;5;187m░\033[38;5;166;48;5;240m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▒\033[38;5;130;48;5;242m▓\033[38;5;82;48;5;242m▓\033[38;5;119;48;5;242m▓\033[38;5;65;48;5;242m▓\033[38;5;65;48;5;241m▓\033[38;5;65;48;5;59m▓\033[38;5;191;48;5;59m▓\033[38;5;221;48;5;59m▓\033[38;5;137;48;5;241m▓\033[38;5;202;48;5;242m▓\033[0m \033[0m \033[0m \033[0m \033[38;5;202;48;5;242m▓\033[38;5;47;48;5;59m▓\033[38;5;50;48;5;187m░\033[38;5;95;48;5;180m▓\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;29;48;5;180m▒\033[38;5;87;48;5;223m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;235m▒\033[38;5;73;48;5;145m▒\033[38;5;51;48;5;230m░\033[38;5;174;48;5;223m▒\033[38;5;221;48;5;223m░\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;84;48;5;180m▒\033[38;5;50;48;5;186m▒\033[38;5;57;48;5;187m▒\033[38;5;51;48;5;187m░\033[38;5;80;48;5;187m░\033[38;5;47;48;5;242m▓\033[38;5;209;48;5;240m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;42;48;5;244m▓\033[38;5;51;48;5;255m░\033[38;5;50;48;5;224m▒\033[38;5;94;48;5;187m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;173m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;179;48;5;180m▒\033[38;5;50;48;5;187m░\033[38;5;29;48;5;242m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;87;48;5;255m░\033[38;5;29;48;5;224m░\033[38;5;172;48;5;223m░\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;143m▒\033[38;5;68;48;5;180m▒\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;248m▒\033[38;5;214;48;5;224m░\033[38;5;214;48;5;186m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;51;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;51;48;5;255m░\033[38;5;220;48;5;187m▒\033[38;5;220;48;5;143m▒\033[38;5;178;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;220;48;5;143m▒\033[38;5;51;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;255m░\033[38;5;172;48;5;187m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;178;48;5;143m▒\033[38;5;80;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;236m▒\033[38;5;69;48;5;223m░\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;172;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;178;48;5;179m▒\033[38;5;42;48;5;179m▒\033[38;5;36;48;5;101m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;230m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;50;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;236m▒\033[38;5;185;48;5;187m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;163;48;5;180m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;235m▒\033[38;5;130;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;32;48;5;179m▒\033[38;5;47;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;224m░\033[38;5;179;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;67;48;5;179m▒\033[38;5;78;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;50;48;5;223m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;25;48;5;179m▒\033[38;5;72;48;5;101m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m▒\033[38;5;179;48;5;223m░\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;67;48;5;180m▒\033[38;5;130;48;5;241m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;230m░\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;50;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;93;48;5;223m░\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;173m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;118;48;5;223m▒\033[38;5;84;48;5;243m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;45;48;5;223m░\033[38;5;136;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;237m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;233m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;235m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;240m▒\033[38;5;94;48;5;101m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;221;48;5;234m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;45;48;5;186m▒\033[38;5;65;48;5;243m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;99;48;5;187m▓\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;52;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;242;48;5;241m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;232;48;5;232m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;252;48;5;252m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;221;48;5;232m \033[38;5;221;48;5;101m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;234;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;238;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;101m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;57;48;5;180m░\033[38;5;113;48;5;243m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;51;48;5;187m░\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;52;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;236;48;5;236m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;234;48;5;234m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;250;48;5;250m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;248;48;5;248m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;236;48;5;236m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;50;48;5;186m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;52;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;245;48;5;245m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;236;48;5;236m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;249;48;5;249m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;241;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;237;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;249;48;5;249m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;50;48;5;223m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;223m░\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;75;48;5;180m░\033[38;5;50;48;5;222m░\033[38;5;35;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;52;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;245;48;5;245m▓\033[38;5;102;48;5;102m▓\033[38;5;102;48;5;102m▓\033[38;5;247;48;5;247m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;235;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;235;48;5;235m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;239;48;5;239m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;242;48;5;241m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;130;48;5;232m \033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;31;48;5;179m░\033[38;5;78;48;5;101m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;50;48;5;187m░\033[0m \033[0m \033[0m \033[38;5;86;48;5;138m▓\033[38;5;50;48;5;186m░\033[38;5;136;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;209;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;237;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;246;48;5;246m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;236;48;5;235m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;232;48;5;232m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;234;48;5;234m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;230;48;5;180m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;230m░\033[38;5;178;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;47;48;5;180m▒\033[38;5;202;48;5;239m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;249m▒\033[38;5;62;48;5;186m░\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;209;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;245;48;5;245m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;234;48;5;234m▓\033[38;5;16;48;5;16m▓\033[38;5;240;48;5;240m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;249;48;5;249m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;251;48;5;251m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;234;48;5;234m▓\033[38;5;233;48;5;233m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;237;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;172;48;5;95m▓\033[38;5;49;48;5;187m▒\033[38;5;208;48;5;223m░\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;179m▒\033[38;5;130;48;5;173m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;42;48;5;95m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;204;48;5;180m▓\033[38;5;220;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;32;48;5;186m▒\033[38;5;87;48;5;229m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;144m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;216;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;234m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;242;48;5;242m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;238;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;232;48;5;232m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;252;48;5;252m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;234;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;50;48;5;187m░\033[38;5;1;48;5;232m░\033[0m \033[38;5;50;48;5;252m▒\033[38;5;190;48;5;187m░\033[38;5;130;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;165;48;5;180m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;223m░\033[38;5;136;48;5;144m▒\033[38;5;178;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;178;48;5;179m▒\033[38;5;50;48;5;187m░\033[38;5;131;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[38;5;51;48;5;223m░\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;233m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;202;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;209;48;5;16m \033[38;5;94;48;5;179m▒\033[38;5;214;48;5;95m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;239m▓\033[38;5;35;48;5;187m░\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[38;5;123;48;5;230m░\033[38;5;26;48;5;186m░\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;200;48;5;180m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;50;48;5;180m░\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;50;48;5;187m░\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;224m░\033[38;5;214;48;5;144m▓\033[38;5;214;48;5;137m▓\033[38;5;94;48;5;233m▒\033[38;5;202;48;5;16m \033[38;5;202;48;5;16m \033[38;5;166;48;5;16m \033[38;5;94;48;5;232m░\033[38;5;94;48;5;137m▓\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;143m▒\033[38;5;94;48;5;233m▒\033[38;5;166;48;5;232m \033[38;5;202;48;5;16m \033[38;5;209;48;5;16m \033[38;5;214;48;5;234m░\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;58m▒\033[38;5;202;48;5;16m \033[38;5;209;48;5;16m \033[38;5;209;48;5;16m \033[38;5;166;48;5;232m \033[38;5;94;48;5;239m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;236m▒\033[38;5;172;48;5;232m \033[38;5;216;48;5;16m \033[38;5;222;48;5;232m \033[38;5;221;48;5;235m▒\033[38;5;221;48;5;95m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;237m▒\033[38;5;222;48;5;233m░\033[38;5;209;48;5;16m \033[38;5;172;48;5;232m \033[38;5;179;48;5;236m▒\033[38;5;214;48;5;101m▓\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;77;48;5;180m▒\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;191;48;5;180m░\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;156;48;5;180m░\033[38;5;84;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;88;48;5;232m░\033[38;5;71;48;5;180m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;51;48;5;223m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;181m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;179;48;5;180m░\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;186m░\033[38;5;178;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;50;48;5;223m░\033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;230m░\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;45;48;5;180m░\033[38;5;84;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;88;48;5;232m░\033[38;5;69;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;47;48;5;186m░\033[38;5;166;48;5;240m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;144m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;179;48;5;180m░\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;221;48;5;222m░\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;167;48;5;232m░\033[0m \033[0m \033[0m \033[38;5;87;48;5;223m░\033[38;5;220;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;80;48;5;180m░\033[38;5;84;48;5;243m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;88;48;5;232m░\033[38;5;29;48;5;180m▓\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;214;48;5;186m▒\033[38;5;50;48;5;224m░\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;93;48;5;186m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m░\033[38;5;178;48;5;186m░\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;87;48;5;230m░\033[0m \033[0m \033[0m \033[38;5;47;48;5;186m▒\033[38;5;221;48;5;143m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;45;48;5;180m░\033[38;5;84;48;5;243m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;50;48;5;181m░\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;186m▒\033[38;5;50;48;5;224m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;186m░\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m░\033[38;5;221;48;5;222m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;50;48;5;223m░\033[0m \033[0m \033[38;5;50;48;5;253m░\033[38;5;214;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;45;48;5;180m▒\033[38;5;84;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;144m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;99;48;5;186m▒\033[38;5;131;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;223m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;50;48;5;223m░\033[0m \033[0m \033[38;5;80;48;5;187m░\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;31;48;5;180m▓\033[38;5;209;48;5;240m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;178;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;87;48;5;229m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;51;48;5;187m░\033[38;5;88;48;5;232m░\033[0m \033[38;5;80;48;5;253m░\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;143m▒\033[38;5;50;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;50;48;5;180m░\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;50;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;223m░\033[38;5;87;48;5;230m░\033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;221;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;144m▒\033[38;5;86;48;5;101m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;88;48;5;232m░\033[38;5;50;48;5;186m░\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;50;48;5;224m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;50;48;5;223m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;99;48;5;180m░\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;206;48;5;180m░\033[38;5;138;48;5;239m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m░\033[38;5;178;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;137m▓\033[38;5;80;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;223m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;185m░\033[38;5;50;48;5;223m░\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;102m▓\033[38;5;178;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;29;48;5;101m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;109;48;5;245m▓\033[38;5;220;48;5;143m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;137m▒\033[38;5;80;48;5;186m░\033[38;5;88;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;252m▒\033[38;5;78;48;5;187m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;50;48;5;223m░\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;95;48;5;240m▓\033[38;5;44;48;5;180m░\033[38;5;221;48;5;137m▓\033[38;5;214;48;5;143m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;220;48;5;180m▒\033[38;5;116;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;50;48;5;144m░\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;143m▒\033[38;5;220;48;5;137m▒\033[38;5;220;48;5;137m▒\033[38;5;220;48;5;137m▒\033[38;5;80;48;5;187m░\033[38;5;88;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;251m▒\033[38;5;214;48;5;180m▒\033[38;5;220;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;52;48;5;180m░\033[38;5;103;48;5;186m▓\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;50;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;186m░\033[38;5;178;48;5;143m▓\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;43;48;5;180m░\033[38;5;43;48;5;102m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;101m▓\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;62;48;5;101m░\033[38;5;29;48;5;243m▓\033[0m \033[0m \033[0m \033[38;5;202;48;5;241m▓\033[38;5;86;48;5;179m▒\033[38;5;220;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;50;48;5;186m░\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[38;5;174;48;5;236m▒\033[38;5;50;48;5;186m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;50;48;5;180m░\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[38;5;209;48;5;239m▓\033[38;5;44;48;5;144m░\033[38;5;178;48;5;143m▓\033[38;5;136;48;5;143m▓\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;187m▒\033[38;5;44;48;5;187m░\033[38;5;138;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▓\033[38;5;161;48;5;187m░\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;220;48;5;143m▒\033[38;5;136;48;5;143m▓\033[38;5;179;48;5;137m▒\033[38;5;130;48;5;137m▓\033[38;5;42;48;5;243m▓\033[0m \033[0m \033[0m \033[38;5;50;48;5;187m▒\033[38;5;220;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;50;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;78;48;5;242m▓\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;69;48;5;179m░\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[38;5;116;48;5;144m▒\033[38;5;136;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;214;48;5;187m▒\033[38;5;50;48;5;250m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;51;48;5;230m░\033[38;5;94;48;5;187m▒\033[38;5;214;48;5;187m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;214;48;5;137m▒\033[38;5;39;48;5;101m▒\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[38;5;80;48;5;187m▒\033[38;5;178;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;114;48;5;179m▒\033[38;5;116;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;186m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;50;48;5;187m░\033[0m \033[0m \033[38;5;116;48;5;249m▒\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;209;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;224m░\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;137m▒\033[38;5;86;48;5;137m▒\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;178;48;5;179m▒\033[38;5;80;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m░\033[38;5;214;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;50;48;5;180m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[38;5;50;48;5;245m▒\033[38;5;214;48;5;101m▓\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;143m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;84;48;5;187m▒\033[38;5;131;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;239m▓\033[38;5;33;48;5;187m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;101m▒\033[38;5;221;48;5;58m▒\033[38;5;94;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;50;48;5;138m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;82;48;5;180m░\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;42;48;5;241m▓\033[38;5;179;48;5;143m▒\033[38;5;214;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;27;48;5;179m░\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[0m \033[38;5;138;48;5;239m▓\033[38;5;85;48;5;137m░\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m░\033[38;5;214;48;5;186m░\033[38;5;214;48;5;186m░\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;47;48;5;187m░\033[38;5;50;48;5;249m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;51;48;5;187m░\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m░\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;186m░\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;144m▓\033[38;5;50;48;5;180m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;180m░\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;50;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;47;48;5;243m▓\033[38;5;57;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;178;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;173m▒\033[38;5;36;48;5;223m░\033[0m \033[0m \033[0m \033[0m \033[38;5;116;48;5;249m▒\033[38;5;136;48;5;95m▓\033[38;5;221;48;5;95m▒\033[38;5;94;48;5;94m▒\033[38;5;214;48;5;101m▒\033[38;5;214;48;5;144m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;186m░\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;199;48;5;187m▒\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;51;48;5;223m░\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;180m▒\033[38;5;136;48;5;187m▒\033[38;5;221;48;5;223m░\033[38;5;221;48;5;187m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;178;48;5;180m▒\033[38;5;221;48;5;144m▓\033[38;5;80;48;5;254m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;138;48;5;238m▓\033[38;5;40;48;5;179m░\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;80;48;5;186m░\033[38;5;131;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;138;48;5;238m▓\033[38;5;200;48;5;186m▓\033[38;5;214;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;208;48;5;180m▓\033[38;5;174;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▓\033[38;5;32;48;5;137m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;178;48;5;222m░\033[38;5;220;48;5;180m▒\033[38;5;220;48;5;180m▒\033[38;5;80;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;246m▓\033[38;5;77;48;5;138m░\033[38;5;136;48;5;144m▓\033[38;5;83;48;5;223m░\033[38;5;136;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;220;48;5;180m▒\033[38;5;69;48;5;180m░\033[38;5;80;48;5;253m░\033[38;5;209;48;5;236m▓\033[38;5;80;48;5;253m░\033[38;5;131;48;5;237m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;84;48;5;180m░\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;137m▒\033[38;5;136;48;5;143m▒\033[38;5;178;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;50;48;5;180m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m░\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;50;48;5;223m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m▒\033[38;5;220;48;5;144m▓\033[38;5;178;48;5;144m▓\033[38;5;221;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;187m▒\033[38;5;94;48;5;186m▒\033[38;5;136;48;5;187m▒\033[38;5;27;48;5;187m░\033[38;5;119;48;5;101m░\033[38;5;116;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;131;48;5;237m▓\033[38;5;131;48;5;237m▓\033[38;5;87;48;5;255m░\033[38;5;87;48;5;254m░\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;50;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;149;48;5;243m▓\033[38;5;101;48;5;187m▓\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;162;48;5;180m▒\033[38;5;174;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▒\033[0m \033[38;5;131;48;5;237m▓\033[38;5;80;48;5;187m░\033[38;5;86;48;5;187m░\033[38;5;220;48;5;187m░\033[38;5;80;48;5;253m░\033[38;5;131;48;5;237m▓\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;185;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;50;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;101;48;5;243m▓\033[38;5;156;48;5;180m░\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;50;48;5;180m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;123;48;5;230m░\033[38;5;214;48;5;143m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;62;48;5;180m░\033[38;5;167;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;137;48;5;243m▓\033[38;5;192;48;5;181m░\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;178;48;5;180m▒\033[38;5;178;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;50;48;5;181m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;214;48;5;143m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;50;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;211;48;5;187m░\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;220;48;5;179m▒\033[38;5;220;48;5;143m▒\033[38;5;50;48;5;187m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;204;48;5;180m░\033[38;5;221;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;69;48;5;143m░\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m░\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;144m▒\033[38;5;87;48;5;224m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;161;48;5;143m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;244m▓\033[38;5;35;48;5;180m░\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;50;48;5;180m░\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;224m░\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;40;48;5;180m░\033[38;5;50;48;5;253m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;45;48;5;241m▓\033[38;5;25;48;5;138m░\033[38;5;179;48;5;137m▓\033[38;5;179;48;5;144m▒\033[38;5;221;48;5;180m▒\033[38;5;178;48;5;180m▒\033[38;5;143;48;5;180m▒\033[38;5;93;48;5;150m▒\033[38;5;80;48;5;187m░\033[38;5;116;48;5;250m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;224m░\033[38;5;178;48;5;144m▓\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;51;48;5;143m░\033[38;5;45;48;5;143m░\033[38;5;80;48;5;143m▒\033[38;5;45;48;5;144m░\033[38;5;50;48;5;145m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;88;48;5;232m░\033[38;5;88;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m");

				$display("\n\033[1;32mCongratulations! Your critical path is below 3!\033[m\n");	
			end
			else begin
		      	$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;246m▓\033[38;5;87;48;5;255m░\033[38;5;87;48;5;230m░\033[38;5;123;48;5;231m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;236m▓\033[38;5;50;48;5;186m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;36;48;5;179m▒\033[38;5;131;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;244m▓\033[38;5;43;48;5;95m▒\033[38;5;50;48;5;186m░\033[38;5;86;48;5;94m░\033[38;5;43;48;5;95m▒\033[38;5;50;48;5;102m▓\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;209;48;5;179m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;172m░\033[38;5;179;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;76;48;5;222m░\033[38;5;66;48;5;247m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;101m▒\033[38;5;156;48;5;173m░\033[38;5;172;48;5;136m░\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;79;48;5;179m▒\033[38;5;73;48;5;248m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;255m░\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;31;48;5;186m░\033[38;5;50;48;5;102m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;138;48;5;239m▓\033[38;5;50;48;5;180m░\033[38;5;172;48;5;136m▒\033[38;5;130;48;5;130m░\033[38;5;172;48;5;130m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;136m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;50;48;5;187m░\033[38;5;50;48;5;244m▓\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;234m▒\033[38;5;90;48;5;179m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;172m░\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;45;48;5;222m░\033[38;5;50;48;5;102m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;202;48;5;235m▓\033[38;5;119;48;5;137m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;172;48;5;130m░\033[38;5;179;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;165;48;5;186m░\033[38;5;109;48;5;246m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▓\033[38;5;50;48;5;144m░\033[38;5;179;48;5;173m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;173m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;38;48;5;186m▒\033[38;5;50;48;5;101m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m▒\033[38;5;50;48;5;143m░\033[38;5;130;48;5;130m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;172;48;5;130m░\033[38;5;172;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;50;48;5;180m░\033[38;5;73;48;5;249m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;238m▓\033[38;5;50;48;5;187m░\033[38;5;179;48;5;173m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;41;48;5;186m░\033[38;5;50;48;5;101m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;50;48;5;187m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;172;48;5;130m░\033[38;5;172;48;5;130m░\033[38;5;172;48;5;130m░\033[38;5;172;48;5;136m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;166;48;5;186m▒\033[38;5;50;48;5;102m▓\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;237m▓\033[38;5;130;48;5;179m▓\033[38;5;179;48;5;172m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;172m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;50;48;5;101m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;173;48;5;179m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;130m░\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;136m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;50;48;5;101m▒\033[38;5;50;48;5;242m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;148;48;5;59m▓\033[38;5;50;48;5;186m░\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;172m░\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;50;48;5;144m▒\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;26;48;5;137m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;130m░\033[38;5;130;48;5;130m░\033[38;5;130;48;5;130m░\033[38;5;172;48;5;130m▒\033[38;5;172;48;5;130m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;101m▒\033[38;5;172;48;5;130m▒\033[38;5;172;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;136m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;80;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;242;48;5;242m▓\033[38;5;50;48;5;186m░\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m░\033[38;5;172;48;5;172m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;172m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;50;48;5;223m░\033[38;5;138;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;231m░\033[38;5;130;48;5;130m░\033[38;5;130;48;5;130m░\033[38;5;172;48;5;130m░\033[38;5;172;48;5;130m░\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;130m▒\033[38;5;172;48;5;101m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;172;48;5;136m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;130m░\033[38;5;179;48;5;136m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;204;48;5;180m▓\033[38;5;109;48;5;247m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;88;48;5;232m░\033[38;5;167;48;5;233m░\033[38;5;167;48;5;233m░\033[38;5;167;48;5;233m░\033[38;5;1;48;5;232m░\033[38;5;1;48;5;232m░\033[38;5;87;48;5;255m░\033[38;5;51;48;5;187m░\033[38;5;50;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;172m▒\033[38;5;172;48;5;172m░\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;50;48;5;223m░\033[38;5;167;48;5;233m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;255m░\033[38;5;172;48;5;130m░\033[38;5;130;48;5;130m░\033[38;5;172;48;5;130m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;101m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;136m▒\033[38;5;179;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;172;48;5;136m▒\033[38;5;130;48;5;94m░\033[38;5;172;48;5;130m░\033[38;5;179;48;5;136m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;136m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;179m▒\033[38;5;185;48;5;180m░\033[38;5;36;48;5;95m▒\033[38;5;42;48;5;238m▓\033[38;5;65;48;5;240m▓\033[38;5;137;48;5;240m▓\033[38;5;202;48;5;59m▓\033[38;5;65;48;5;240m▓\033[38;5;72;48;5;238m▓\033[38;5;50;48;5;181m▒\033[38;5;50;48;5;223m░\033[38;5;50;48;5;223m░\033[38;5;50;48;5;223m░\033[38;5;50;48;5;223m░\033[38;5;50;48;5;186m░\033[38;5;50;48;5;186m░\033[38;5;205;48;5;186m░\033[38;5;167;48;5;186m▒\033[38;5;38;48;5;180m▒\033[38;5;48;48;5;179m▒\033[38;5;114;48;5;179m▒\033[38;5;114;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;38;48;5;186m▓\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;254m░\033[38;5;130;48;5;130m░\033[38;5;172;48;5;130m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;130m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;130m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;130m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;172;48;5;130m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;136m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;173m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;116;48;5;249m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;255m░\033[38;5;130;48;5;130m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;130m░\033[38;5;172;48;5;130m░\033[38;5;172;48;5;136m░\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;172;48;5;235m▒\033[38;5;130;48;5;58m▒\033[38;5;208;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;130m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;136m▒\033[38;5;172;48;5;136m▒\033[38;5;130;48;5;130m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;130;48;5;130m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;172m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;51;48;5;187m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;109;48;5;247m▓\033[38;5;172;48;5;130m░\033[38;5;130;48;5;130m░\033[38;5;130;48;5;130m░\033[38;5;172;48;5;130m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;236m▒\033[38;5;130;48;5;236m░\033[38;5;130;48;5;236m░\033[38;5;130;48;5;235m▒\033[38;5;172;48;5;235m▒\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;172;48;5;130m▒\033[38;5;172;48;5;136m░\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;172;48;5;136m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;130;48;5;130m░\033[38;5;172;48;5;130m░\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;215m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;50;48;5;223m░\033[38;5;116;48;5;250m▒\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;99;48;5;137m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;130m░\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;236m▒\033[38;5;172;48;5;236m░\033[38;5;172;48;5;234m▒\033[38;5;172;48;5;234m▒\033[38;5;130;48;5;235m▒\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;136m▒\033[38;5;172;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;136m▒\033[38;5;130;48;5;130m░\033[38;5;130;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;221m░\033[38;5;94;48;5;221m░\033[38;5;94;48;5;185m░\033[38;5;68;48;5;186m▒\033[38;5;50;48;5;144m▒\033[38;5;73;48;5;247m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;209;48;5;180m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;236m▒\033[38;5;172;48;5;235m▒\033[38;5;214;48;5;233m▒\033[38;5;221;48;5;233m░\033[38;5;220;48;5;234m▒\033[38;5;172;48;5;238m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;136m▒\033[38;5;130;48;5;130m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;172;48;5;136m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;136m░\033[38;5;179;48;5;172m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;215m░\033[38;5;214;48;5;179m░\033[38;5;43;48;5;186m▒\033[38;5;51;48;5;230m░\033[38;5;109;48;5;245m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;87;48;5;224m░\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;136m░\033[38;5;179;48;5;136m░\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;236m▒\033[38;5;172;48;5;236m▒\033[38;5;130;48;5;235m▒\033[38;5;179;48;5;234m▒\033[38;5;94;48;5;233m░\033[38;5;221;48;5;233m░\033[38;5;94;48;5;235m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;130m▒\033[38;5;172;48;5;130m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;130m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;172m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;222m░\033[38;5;221;48;5;186m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;186m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;186m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;221m░\033[38;5;94;48;5;185m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;221m░\033[38;5;161;48;5;222m░\033[38;5;51;48;5;230m░\033[38;5;166;48;5;236m▓\033[38;5;209;48;5;237m▓\033[38;5;174;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;235m▒\033[38;5;50;48;5;187m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;214;48;5;136m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;236m▒\033[38;5;130;48;5;235m▒\033[38;5;172;48;5;234m▒\033[38;5;179;48;5;234m▒\033[38;5;221;48;5;233m░\033[38;5;221;48;5;233m░\033[38;5;172;48;5;234m░\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;136m▒\033[38;5;130;48;5;130m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;136m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;172m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;172m░\033[38;5;179;48;5;136m░\033[38;5;179;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;198;48;5;222m▒\033[38;5;116;48;5;249m▒\033[38;5;88;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;235m▒\033[38;5;50;48;5;187m░\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;136m░\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;94;48;5;173m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;172;48;5;136m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;239m▒\033[38;5;179;48;5;235m▒\033[38;5;172;48;5;235m▒\033[38;5;214;48;5;234m▒\033[38;5;214;48;5;234m▒\033[38;5;214;48;5;234m▒\033[38;5;94;48;5;234m▒\033[38;5;179;48;5;234m▒\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;95m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;172m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;172m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;136m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;222m░\033[38;5;94;48;5;186m░\033[38;5;221;48;5;222m░\033[38;5;221;48;5;186m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;50;48;5;223m░\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m▒\033[38;5;78;48;5;179m▒\033[38;5;172;48;5;136m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;136m▒\033[38;5;130;48;5;130m░\033[38;5;172;48;5;130m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;235m▒\033[38;5;130;48;5;58m░\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;173m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;172m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;221m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;50;48;5;223m░\033[38;5;174;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;87;48;5;230m░\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;94;48;5;137m▒\033[38;5;172;48;5;95m▒\033[38;5;130;48;5;58m▒\033[38;5;130;48;5;94m░\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m░\033[38;5;179;48;5;136m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;130m░\033[38;5;130;48;5;130m░\033[38;5;172;48;5;130m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;136m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;173m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;173m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;221m░\033[38;5;165;48;5;186m▒\033[38;5;95;48;5;241m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;223m░\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;136m▒\033[38;5;172;48;5;136m░\033[38;5;179;48;5;136m▒\033[38;5;172;48;5;136m░\033[38;5;179;48;5;136m░\033[38;5;179;48;5;136m░\033[38;5;179;48;5;136m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;136m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;137m▒\033[38;5;172;48;5;136m░\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m░\033[38;5;179;48;5;172m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;178;48;5;144m▓\033[38;5;178;48;5;101m▓\033[38;5;94;48;5;240m▓\033[38;5;179;48;5;239m▒\033[38;5;130;48;5;94m▒\033[38;5;179;48;5;240m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;221m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;116;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;162;48;5;180m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;172;48;5;172m▒\033[38;5;172;48;5;130m░\033[38;5;172;48;5;130m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;172;48;5;130m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;136m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;143m▓\033[38;5;136;48;5;101m▓\033[38;5;221;48;5;236m▒\033[38;5;136;48;5;232m \033[38;5;222;48;5;16m \033[38;5;221;48;5;16m \033[38;5;136;48;5;232m \033[38;5;136;48;5;233m▒\033[38;5;178;48;5;233m▒\033[38;5;136;48;5;234m▒\033[38;5;221;48;5;137m▓\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;185m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;50;48;5;144m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;144m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;172m░\033[38;5;172;48;5;136m░\033[38;5;130;48;5;130m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;130m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;172m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;136m▒\033[38;5;214;48;5;136m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;95m▒\033[38;5;179;48;5;236m▒\033[38;5;136;48;5;237m▓\033[38;5;178;48;5;246m▓\033[38;5;221;48;5;232m \033[38;5;94;48;5;235m▒\033[38;5;221;48;5;240m▓\033[38;5;178;48;5;101m▓\033[38;5;221;48;5;239m▓\033[38;5;220;48;5;144m▓\033[38;5;221;48;5;95m▓\033[38;5;136;48;5;143m▓\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;222m░\033[38;5;136;48;5;223m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;229m░\033[38;5;178;48;5;223m░\033[38;5;221;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;99;48;5;223m▒\033[38;5;66;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;137m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;172m▒\033[38;5;172;48;5;136m░\033[38;5;130;48;5;130m░\033[38;5;130;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;130m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;101m▒\033[38;5;221;48;5;137m▓\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;236m▒\033[38;5;94;48;5;232m░\033[38;5;178;48;5;232m \033[38;5;221;48;5;232m░\033[38;5;94;48;5;233m░\033[38;5;179;48;5;235m▒\033[38;5;179;48;5;235m▒\033[38;5;221;48;5;233m▒\033[38;5;94;48;5;237m▓\033[38;5;220;48;5;187m▒\033[38;5;136;48;5;101m▓\033[38;5;178;48;5;180m▓\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m \033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m \033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;136;48;5;223m░\033[38;5;221;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;50;48;5;187m░\033[38;5;138;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;244m▓\033[38;5;78;48;5;186m▓\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;172m░\033[38;5;172;48;5;136m░\033[38;5;130;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;172;48;5;130m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;101m▒\033[38;5;214;48;5;239m▓\033[38;5;221;48;5;234m▒\033[38;5;136;48;5;232m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;220;48;5;232m \033[38;5;221;48;5;232m \033[38;5;136;48;5;235m▒\033[38;5;136;48;5;95m▓\033[38;5;136;48;5;137m▓\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;136;48;5;233m░\033[38;5;222;48;5;16m \033[38;5;221;48;5;232m \033[38;5;221;48;5;234m▒\033[38;5;94;48;5;237m▒\033[38;5;94;48;5;237m▓\033[38;5;214;48;5;236m▒\033[38;5;136;48;5;241m▓\033[38;5;220;48;5;144m▓\033[38;5;221;48;5;95m▓\033[38;5;178;48;5;144m▓\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;220;48;5;230m░\033[38;5;178;48;5;229m░\033[38;5;221;48;5;223m░\033[38;5;21;48;5;223m░\033[38;5;29;48;5;239m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;50;48;5;137m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;172m░\033[38;5;172;48;5;136m░\033[38;5;130;48;5;130m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;172;48;5;130m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;172m▒\033[38;5;172;48;5;136m▒\033[38;5;179;48;5;137m▒\033[38;5;94;48;5;101m▒\033[38;5;221;48;5;237m▒\033[38;5;130;48;5;16m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;136;48;5;232m \033[38;5;136;48;5;233m▒\033[38;5;178;48;5;238m▓\033[38;5;220;48;5;248m▓\033[38;5;220;48;5;187m▓\033[38;5;220;48;5;144m▓\033[38;5;221;48;5;240m▓\033[38;5;220;48;5;235m▓\033[38;5;220;48;5;234m▒\033[38;5;214;48;5;239m▒\033[38;5;94;48;5;101m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;238m▒\033[38;5;214;48;5;234m▒\033[38;5;94;48;5;236m▒\033[38;5;94;48;5;236m▒\033[38;5;214;48;5;235m▒\033[38;5;136;48;5;235m▒\033[38;5;221;48;5;95m▓\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;144m▓\033[38;5;178;48;5;186m▒\033[38;5;221;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;136;48;5;223m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m \033[38;5;220;48;5;230m \033[38;5;230;48;5;230m \033[38;5;220;48;5;230m░\033[38;5;220;48;5;229m░\033[38;5;136;48;5;223m░\033[38;5;221;48;5;222m░\033[38;5;51;48;5;230m░\033[38;5;131;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;101;48;5;239m▓\033[38;5;60;48;5;186m▓\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;172m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;130m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;130m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;130m▒\033[38;5;179;48;5;58m▒\033[38;5;215;48;5;232m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;221;48;5;232m░\033[38;5;136;48;5;232m \033[38;5;215;48;5;16m \033[38;5;221;48;5;16m \033[38;5;136;48;5;232m \033[38;5;221;48;5;233m░\033[38;5;221;48;5;233m░\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;181m▓\033[38;5;178;48;5;144m▓\033[38;5;220;48;5;237m▓\033[38;5;172;48;5;16m \033[38;5;221;48;5;233m░\033[38;5;179;48;5;235m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;136m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;186m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;186m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;179;48;5;215m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;221m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;240m▒\033[38;5;179;48;5;95m▓\033[38;5;136;48;5;101m▓\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;220;48;5;230m \033[38;5;220;48;5;230m░\033[38;5;220;48;5;229m░\033[38;5;99;48;5;223m▒\033[38;5;131;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;42;48;5;238m▓\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;101m▒\033[38;5;172;48;5;236m▒\033[38;5;214;48;5;235m▒\033[38;5;220;48;5;233m░\033[38;5;94;48;5;232m░\033[38;5;94;48;5;232m \033[38;5;222;48;5;232m \033[38;5;178;48;5;16m \033[38;5;215;48;5;16m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;215;48;5;16m \033[38;5;136;48;5;237m▓\033[38;5;178;48;5;137m▓\033[38;5;136;48;5;144m▓\033[38;5;178;48;5;101m▓\033[38;5;136;48;5;234m▒\033[38;5;222;48;5;16m \033[38;5;136;48;5;233m░\033[38;5;179;48;5;234m▒\033[38;5;130;48;5;58m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;172;48;5;136m░\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;185m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;185m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;186m░\033[38;5;178;48;5;223m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m \033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m \033[38;5;220;48;5;230m░\033[38;5;220;48;5;229m░\033[38;5;178;48;5;223m░\033[38;5;87;48;5;230m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;236m▒\033[38;5;50;48;5;223m░\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;59m▓\033[38;5;221;48;5;239m▓\033[38;5;136;48;5;239m▓\033[38;5;220;48;5;232m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;94;48;5;232m \033[38;5;179;48;5;233m░\033[38;5;214;48;5;235m▒\033[38;5;179;48;5;234m▒\033[38;5;221;48;5;237m▓\033[38;5;94;48;5;95m▓\033[38;5;136;48;5;101m▓\033[38;5;94;48;5;237m▓\033[38;5;221;48;5;233m░\033[38;5;94;48;5;236m▒\033[38;5;179;48;5;234m▒\033[38;5;172;48;5;58m▒\033[38;5;214;48;5;101m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;186m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;221m░\033[38;5;179;48;5;215m░\033[38;5;214;48;5;215m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;222m░\033[38;5;94;48;5;186m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;221;48;5;222m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;229m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m \033[38;5;220;48;5;230m \033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m \033[38;5;220;48;5;230m░\033[38;5;220;48;5;229m░\033[38;5;178;48;5;223m░\033[38;5;87;48;5;231m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;236m▒\033[38;5;50;48;5;187m░\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;144m▓\033[38;5;136;48;5;101m▓\033[38;5;221;48;5;59m▓\033[38;5;221;48;5;238m▓\033[38;5;221;48;5;238m▓\033[38;5;221;48;5;239m▓\033[38;5;178;48;5;240m▓\033[38;5;136;48;5;238m▓\033[38;5;94;48;5;237m▓\033[38;5;221;48;5;95m▓\033[38;5;221;48;5;240m▓\033[38;5;214;48;5;236m▒\033[38;5;172;48;5;234m▒\033[38;5;94;48;5;236m▒\033[38;5;221;48;5;95m▓\033[38;5;179;48;5;95m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;136m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;214;48;5;221m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;214;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;229m░\033[38;5;215;48;5;230m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;236m▒\033[38;5;170;48;5;186m░\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;143m▓\033[38;5;221;48;5;143m▓\033[38;5;136;48;5;143m▓\033[38;5;221;48;5;137m▓\033[38;5;221;48;5;137m▓\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;186m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;222m░\033[38;5;136;48;5;223m░\033[38;5;221;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;136;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;41;48;5;230m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;235m▒\033[38;5;168;48;5;186m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;221;48;5;222m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;222m░\033[38;5;221;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;144m▒\033[38;5;178;48;5;144m▓\033[38;5;136;48;5;144m▓\033[38;5;136;48;5;143m▓\033[38;5;136;48;5;137m▓\033[38;5;136;48;5;144m▓\033[38;5;136;48;5;144m▓\033[38;5;178;48;5;144m▓\033[38;5;220;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m \033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m \033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;229m░\033[38;5;87;48;5;255m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;247m▓\033[38;5;220;48;5;222m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;187m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;136;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;180m▒\033[38;5;178;48;5;180m▓\033[38;5;178;48;5;144m▓\033[38;5;136;48;5;101m▓\033[38;5;221;48;5;240m▓\033[38;5;94;48;5;239m▓\033[38;5;221;48;5;240m▓\033[38;5;221;48;5;240m▓\033[38;5;221;48;5;240m▓\033[38;5;221;48;5;59m▓\033[38;5;221;48;5;95m▓\033[38;5;221;48;5;95m▓\033[38;5;221;48;5;241m▓\033[38;5;221;48;5;59m▓\033[38;5;221;48;5;240m▓\033[38;5;221;48;5;95m▓\033[38;5;136;48;5;101m▓\033[38;5;221;48;5;101m▓\033[38;5;136;48;5;138m▓\033[38;5;220;48;5;187m▓\033[38;5;220;48;5;230m \033[38;5;220;48;5;230m░\033[38;5;220;48;5;229m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;229m░\033[38;5;178;48;5;223m░\033[38;5;80;48;5;249m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;136;48;5;187m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;220;48;5;180m▓\033[38;5;178;48;5;144m▓\033[38;5;221;48;5;95m▓\033[38;5;94;48;5;238m▓\033[38;5;94;48;5;236m▒\033[38;5;179;48;5;235m▒\033[38;5;179;48;5;235m▒\033[38;5;179;48;5;236m▒\033[38;5;214;48;5;235m▒\033[38;5;136;48;5;236m▓\033[38;5;221;48;5;234m▒\033[38;5;221;48;5;233m▒\033[38;5;221;48;5;232m░\033[38;5;136;48;5;232m░\033[38;5;136;48;5;232m \033[38;5;221;48;5;233m░\033[38;5;178;48;5;232m \033[38;5;221;48;5;233m░\033[38;5;94;48;5;232m░\033[38;5;214;48;5;234m▒\033[38;5;94;48;5;234m▒\033[38;5;178;48;5;101m▓\033[38;5;220;48;5;230m▒\033[38;5;220;48;5;230m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;178;48;5;223m░\033[38;5;70;48;5;187m░\033[38;5;50;48;5;245m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;255m░\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;186m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;220;48;5;223m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;94;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;136;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;138m▓\033[38;5;214;48;5;235m▒\033[38;5;214;48;5;235m▒\033[38;5;179;48;5;235m▒\033[38;5;214;48;5;233m▒\033[38;5;221;48;5;232m \033[38;5;222;48;5;16m \033[38;5;130;48;5;16m \033[38;5;130;48;5;232m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;215;48;5;16m \033[38;5;178;48;5;16m \033[38;5;221;48;5;16m \033[38;5;221;48;5;232m \033[38;5;172;48;5;16m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;221;48;5;232m \033[38;5;136;48;5;238m▓\033[38;5;220;48;5;187m▓\033[38;5;220;48;5;230m \033[38;5;220;48;5;230m \033[38;5;220;48;5;230m░\033[38;5;220;48;5;229m░\033[38;5;178;48;5;223m░\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;223m░\033[38;5;220;48;5;229m░\033[38;5;69;48;5;223m▒\033[38;5;116;48;5;245m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;113;48;5;241m▓\033[38;5;35;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;187m▒\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;220;48;5;181m▓\033[38;5;178;48;5;101m▓\033[38;5;221;48;5;237m▓\033[38;5;94;48;5;234m▒\033[38;5;221;48;5;233m░\033[38;5;178;48;5;16m \033[38;5;215;48;5;16m \033[38;5;172;48;5;232m \033[38;5;222;48;5;16m \033[38;5;215;48;5;16m \033[38;5;222;48;5;16m \033[38;5;215;48;5;16m \033[38;5;222;48;5;16m \033[38;5;215;48;5;16m \033[38;5;222;48;5;16m \033[38;5;215;48;5;16m \033[38;5;172;48;5;232m \033[38;5;214;48;5;233m░\033[38;5;178;48;5;16m \033[38;5;215;48;5;16m \033[38;5;220;48;5;232m \033[38;5;136;48;5;235m▒\033[38;5;136;48;5;101m▓\033[38;5;220;48;5;187m▒\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m \033[38;5;178;48;5;223m░\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;220;48;5;187m▒\033[38;5;178;48;5;223m▒\033[38;5;220;48;5;187m▒\033[38;5;80;48;5;181m░\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;245m▓\033[38;5;220;48;5;186m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;187m▓\033[38;5;220;48;5;249m▓\033[38;5;178;48;5;101m▓\033[38;5;221;48;5;238m▓\033[38;5;214;48;5;233m░\033[38;5;221;48;5;16m \033[38;5;222;48;5;16m \033[38;5;130;48;5;16m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;172;48;5;232m \033[38;5;221;48;5;233m░\033[38;5;179;48;5;233m░\033[38;5;221;48;5;232m░\033[38;5;94;48;5;235m▒\033[38;5;221;48;5;238m▓\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;144m▓\033[38;5;178;48;5;101m▓\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;220;48;5;229m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;136;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;230m░\033[38;5;220;48;5;230m░\033[38;5;214;48;5;230m▓\033[38;5;66;48;5;242m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;101m▒\033[38;5;46;48;5;180m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;136m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;220;48;5;187m▓\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;187m▓\033[38;5;220;48;5;187m▓\033[38;5;220;48;5;187m▒\033[38;5;220;48;5;249m▓\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;221;48;5;241m▓\033[38;5;94;48;5;237m▓\033[38;5;214;48;5;235m▒\033[38;5;178;48;5;232m \033[38;5;221;48;5;16m \033[38;5;215;48;5;16m \033[38;5;178;48;5;232m \033[38;5;94;48;5;233m▒\033[38;5;214;48;5;233m░\033[38;5;172;48;5;232m \033[38;5;172;48;5;16m \033[38;5;178;48;5;16m \033[38;5;214;48;5;233m░\033[38;5;178;48;5;232m \033[38;5;221;48;5;16m \033[38;5;221;48;5;232m░\033[38;5;214;48;5;234m▒\033[38;5;94;48;5;233m▒\033[38;5;214;48;5;234m▒\033[38;5;94;48;5;233m▒\033[38;5;136;48;5;240m▓\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;181m▓\033[38;5;220;48;5;187m▓\033[38;5;220;48;5;187m▒\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;51;48;5;230m░\033[38;5;131;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[38;5;36;48;5;242m▓\033[38;5;142;48;5;186m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m░\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;136m▒\033[38;5;214;48;5;136m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;144m▒\033[38;5;178;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;178;48;5;180m▒\033[38;5;178;48;5;144m▓\033[38;5;178;48;5;101m▓\033[38;5;136;48;5;138m▓\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;249m▓\033[38;5;220;48;5;144m▓\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;95m▓\033[38;5;221;48;5;238m▓\033[38;5;214;48;5;237m▓\033[38;5;179;48;5;234m▒\033[38;5;172;48;5;16m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;94;48;5;232m░\033[38;5;94;48;5;233m░\033[38;5;136;48;5;233m░\033[38;5;221;48;5;232m \033[38;5;94;48;5;232m \033[38;5;221;48;5;233m░\033[38;5;221;48;5;233m░\033[38;5;94;48;5;233m▒\033[38;5;94;48;5;235m▒\033[38;5;94;48;5;240m▓\033[38;5;136;48;5;101m▓\033[38;5;178;48;5;144m▓\033[38;5;220;48;5;249m▓\033[38;5;220;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;223m░\033[38;5;51;48;5;230m░\033[38;5;138;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[38;5;138;48;5;237m▓\033[38;5;221;48;5;223m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;172m▒\033[38;5;214;48;5;136m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;187m▓\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;220;48;5;180m▓\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;220;48;5;180m▓\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;178;48;5;144m▓\033[38;5;178;48;5;101m▓\033[38;5;178;48;5;101m▓\033[38;5;136;48;5;101m▓\033[38;5;94;48;5;239m▓\033[38;5;214;48;5;236m▒\033[38;5;214;48;5;237m▓\033[38;5;94;48;5;236m▒\033[38;5;179;48;5;234m▒\033[38;5;221;48;5;233m░\033[38;5;136;48;5;232m \033[38;5;222;48;5;16m \033[38;5;94;48;5;232m \033[38;5;221;48;5;232m \033[38;5;94;48;5;232m \033[38;5;94;48;5;232m \033[38;5;94;48;5;233m▒\033[38;5;214;48;5;234m▒\033[38;5;94;48;5;236m▒\033[38;5;221;48;5;239m▓\033[38;5;221;48;5;95m▓\033[38;5;136;48;5;101m▓\033[38;5;178;48;5;101m▓\033[38;5;178;48;5;138m▓\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;181m▓\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;223m░\033[38;5;220;48;5;223m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;223m░\033[38;5;136;48;5;187m▒\033[38;5;51;48;5;224m░\033[38;5;138;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[38;5;41;48;5;238m▓\033[38;5;80;48;5;186m▒\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;136m▒\033[38;5;214;48;5;136m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;144m▒\033[38;5;136;48;5;180m▒\033[38;5;178;48;5;144m▓\033[38;5;136;48;5;144m▓\033[38;5;178;48;5;144m▓\033[38;5;178;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;249m▓\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;137m▓\033[38;5;221;48;5;95m▓\033[38;5;221;48;5;59m▓\033[38;5;94;48;5;239m▓\033[38;5;94;48;5;236m▒\033[38;5;94;48;5;236m▒\033[38;5;94;48;5;234m▒\033[38;5;179;48;5;234m▒\033[38;5;179;48;5;234m▒\033[38;5;136;48;5;233m░\033[38;5;94;48;5;233m▒\033[38;5;136;48;5;233m░\033[38;5;136;48;5;233m░\033[38;5;94;48;5;234m▒\033[38;5;214;48;5;235m▒\033[38;5;214;48;5;237m▓\033[38;5;94;48;5;238m▓\033[38;5;94;48;5;238m▓\033[38;5;221;48;5;238m▓\033[38;5;136;48;5;59m▓\033[38;5;136;48;5;101m▓\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;223m░\033[38;5;220;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;178;48;5;223m░\033[38;5;51;48;5;230m░\033[38;5;138;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[38;5;167;48;5;233m░\033[38;5;179;48;5;223m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;178;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;178;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;144m▒\033[38;5;136;48;5;144m▒\033[38;5;136;48;5;137m▓\033[38;5;178;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;101m▓\033[38;5;178;48;5;137m▓\033[38;5;221;48;5;240m▓\033[38;5;221;48;5;95m▓\033[38;5;221;48;5;95m▓\033[38;5;214;48;5;236m▒\033[38;5;214;48;5;237m▓\033[38;5;214;48;5;236m▒\033[38;5;179;48;5;235m▒\033[38;5;179;48;5;234m▒\033[38;5;179;48;5;235m▒\033[38;5;94;48;5;237m▓\033[38;5;221;48;5;236m▒\033[38;5;94;48;5;236m▒\033[38;5;94;48;5;236m▒\033[38;5;214;48;5;236m▒\033[38;5;94;48;5;237m▓\033[38;5;94;48;5;237m▓\033[38;5;94;48;5;239m▓\033[38;5;221;48;5;239m▓\033[38;5;94;48;5;239m▓\033[38;5;221;48;5;95m▓\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;137m▓\033[38;5;136;48;5;180m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;220;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;51;48;5;230m░\033[38;5;138;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[38;5;167;48;5;233m▒\033[38;5;106;48;5;223m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;136m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;136m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;144m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;137m▓\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;180m▒\033[38;5;178;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;136;48;5;101m▓\033[38;5;178;48;5;138m▓\033[38;5;221;48;5;95m▓\033[38;5;221;48;5;240m▓\033[38;5;94;48;5;238m▓\033[38;5;94;48;5;236m▒\033[38;5;214;48;5;236m▒\033[38;5;94;48;5;237m▓\033[38;5;94;48;5;238m▓\033[38;5;94;48;5;237m▓\033[38;5;94;48;5;238m▓\033[38;5;94;48;5;237m▓\033[38;5;136;48;5;236m▓\033[38;5;214;48;5;235m▒\033[38;5;94;48;5;236m▒\033[38;5;94;48;5;237m▓\033[38;5;94;48;5;239m▓\033[38;5;221;48;5;239m▓\033[38;5;94;48;5;239m▓\033[38;5;221;48;5;95m▓\033[38;5;94;48;5;59m▓\033[38;5;221;48;5;101m▓\033[38;5;136;48;5;144m▓\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;220;48;5;229m░\033[38;5;178;48;5;229m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;51;48;5;230m░\033[38;5;138;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[38;5;167;48;5;234m▒\033[38;5;51;48;5;223m░\033[38;5;94;48;5;179m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;173m▒\033[38;5;94;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;137m▓\033[38;5;221;48;5;137m▓\033[38;5;136;48;5;137m▓\033[38;5;221;48;5;101m▓\033[38;5;94;48;5;95m▓\033[38;5;221;48;5;59m▓\033[38;5;94;48;5;237m▓\033[38;5;179;48;5;235m▒\033[38;5;94;48;5;238m▓\033[38;5;94;48;5;238m▓\033[38;5;221;48;5;235m▒\033[38;5;221;48;5;237m▓\033[38;5;178;48;5;232m░\033[38;5;222;48;5;16m \033[38;5;215;48;5;16m \033[38;5;222;48;5;16m \033[38;5;215;48;5;16m \033[38;5;222;48;5;16m \033[38;5;221;48;5;16m \033[38;5;221;48;5;233m░\033[38;5;94;48;5;235m▒\033[38;5;94;48;5;237m▓\033[38;5;94;48;5;238m▓\033[38;5;221;48;5;101m▓\033[38;5;178;48;5;180m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;51;48;5;254m░\033[38;5;131;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[38;5;167;48;5;234m▒\033[38;5;51;48;5;224m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▓\033[38;5;221;48;5;137m▓\033[38;5;221;48;5;101m▓\033[38;5;221;48;5;101m▓\033[38;5;221;48;5;101m▓\033[38;5;221;48;5;137m▓\033[38;5;136;48;5;143m▓\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▓\033[38;5;136;48;5;143m▓\033[38;5;136;48;5;143m▓\033[38;5;214;48;5;101m▓\033[38;5;214;48;5;95m▓\033[38;5;94;48;5;239m▓\033[38;5;221;48;5;235m▒\033[38;5;94;48;5;232m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;222;48;5;16m \033[38;5;215;48;5;16m \033[38;5;172;48;5;16m \033[38;5;130;48;5;16m \033[38;5;172;48;5;16m \033[38;5;178;48;5;232m \033[38;5;136;48;5;232m░\033[38;5;221;48;5;233m░\033[38;5;214;48;5;234m▒\033[38;5;179;48;5;235m▒\033[38;5;179;48;5;235m▒\033[38;5;214;48;5;236m▒\033[38;5;94;48;5;237m▓\033[38;5;179;48;5;238m▓\033[38;5;221;48;5;101m▓\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;223m░\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;50;48;5;59m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[38;5;167;48;5;234m▒\033[38;5;87;48;5;230m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;136m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;180m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▓\033[38;5;221;48;5;101m▓\033[38;5;179;48;5;240m▒\033[38;5;94;48;5;236m▒\033[38;5;179;48;5;234m▒\033[38;5;221;48;5;232m \033[38;5;94;48;5;236m▓\033[38;5;221;48;5;233m░\033[38;5;94;48;5;232m \033[38;5;94;48;5;235m▒\033[38;5;214;48;5;236m▒\033[38;5;221;48;5;238m▓\033[38;5;94;48;5;238m▓\033[38;5;94;48;5;95m▓\033[38;5;221;48;5;101m▓\033[38;5;179;48;5;95m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;137m▓\033[38;5;221;48;5;101m▓\033[38;5;94;48;5;237m▓\033[38;5;179;48;5;239m▓\033[38;5;94;48;5;236m▒\033[38;5;221;48;5;232m \033[38;5;136;48;5;232m \033[38;5;221;48;5;232m \033[38;5;130;48;5;16m \033[38;5;94;48;5;233m░\033[38;5;136;48;5;232m \033[38;5;221;48;5;233m░\033[38;5;214;48;5;235m▒\033[38;5;179;48;5;234m▒\033[38;5;214;48;5;233m▒\033[38;5;214;48;5;234m▒\033[38;5;94;48;5;233m▒\033[38;5;179;48;5;234m▒\033[38;5;214;48;5;234m▒\033[38;5;214;48;5;235m▒\033[38;5;94;48;5;236m▒\033[38;5;94;48;5;237m▓\033[38;5;94;48;5;237m▓\033[38;5;94;48;5;240m▓\033[38;5;136;48;5;137m▓\033[38;5;178;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;220;48;5;223m░\033[38;5;105;48;5;230m░\033[38;5;66;48;5;242m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[38;5;137;48;5;235m▓\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;179;48;5;173m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;172m▒\033[38;5;214;48;5;136m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;136m░\033[38;5;214;48;5;136m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;178;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;101m▓\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;179;48;5;240m▓\033[38;5;136;48;5;59m▓\033[38;5;221;48;5;238m▓\033[38;5;94;48;5;235m▒\033[38;5;94;48;5;233m▒\033[38;5;221;48;5;234m▒\033[38;5;179;48;5;234m▒\033[38;5;179;48;5;235m▒\033[38;5;179;48;5;234m▒\033[38;5;172;48;5;234m▒\033[38;5;179;48;5;235m▒\033[38;5;94;48;5;233m▒\033[38;5;214;48;5;233m░\033[38;5;172;48;5;232m \033[38;5;214;48;5;233m░\033[38;5;136;48;5;233m░\033[38;5;214;48;5;235m▒\033[38;5;179;48;5;234m▒\033[38;5;214;48;5;236m▒\033[38;5;214;48;5;236m▒\033[38;5;179;48;5;234m▒\033[38;5;179;48;5;234m▒\033[38;5;179;48;5;234m▒\033[38;5;214;48;5;235m▒\033[38;5;214;48;5;236m▒\033[38;5;94;48;5;234m▒\033[38;5;221;48;5;232m \033[38;5;179;48;5;236m▒\033[38;5;179;48;5;235m▒\033[38;5;214;48;5;236m▒\033[38;5;94;48;5;238m▓\033[38;5;94;48;5;240m▓\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;137m▓\033[38;5;136;48;5;144m▓\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;136;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;81;48;5;229m░\033[38;5;116;48;5;246m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[38;5;209;48;5;237m▓\033[38;5;204;48;5;186m░\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;179;48;5;172m▒\033[38;5;214;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;214;48;5;136m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;95m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;239m▒\033[38;5;172;48;5;58m▒\033[38;5;94;48;5;239m▓\033[38;5;179;48;5;238m▒\033[38;5;94;48;5;237m▒\033[38;5;179;48;5;235m▒\033[38;5;214;48;5;235m▒\033[38;5;214;48;5;235m▒\033[38;5;94;48;5;237m▓\033[38;5;94;48;5;238m▓\033[38;5;221;48;5;238m▓\033[38;5;221;48;5;239m▓\033[38;5;221;48;5;240m▓\033[38;5;94;48;5;238m▓\033[38;5;221;48;5;240m▓\033[38;5;94;48;5;239m▓\033[38;5;214;48;5;239m▓\033[38;5;221;48;5;239m▓\033[38;5;94;48;5;238m▓\033[38;5;172;48;5;238m▒\033[38;5;94;48;5;239m▓\033[38;5;94;48;5;239m▓\033[38;5;214;48;5;240m▓\033[38;5;94;48;5;101m▓\033[38;5;221;48;5;137m▓\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;223m░\033[38;5;136;48;5;187m▒\033[38;5;136;48;5;223m░\033[38;5;136;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;136;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;44;48;5;144m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[38;5;167;48;5;233m▒\033[38;5;221;48;5;101m░\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;136m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;136m▒\033[38;5;172;48;5;136m░\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m░\033[38;5;214;48;5;136m▒\033[38;5;179;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;179;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;101m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;101m▒\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;179;48;5;95m▒\033[38;5;214;48;5;95m▓\033[38;5;221;48;5;101m▓\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;136;48;5;101m▓\033[38;5;179;48;5;101m▒\033[38;5;214;48;5;101m▓\033[38;5;214;48;5;101m▒\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;101m▓\033[38;5;179;48;5;101m▒\033[38;5;221;48;5;59m▓\033[38;5;179;48;5;95m▓\033[38;5;94;48;5;95m▓\033[38;5;94;48;5;101m▓\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;136;48;5;223m░\033[38;5;136;48;5;223m░\033[38;5;221;48;5;223m░\033[38;5;51;48;5;224m░\033[38;5;131;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;247m▓\033[38;5;134;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;173m▒\033[38;5;214;48;5;136m▒\033[38;5;179;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;173m▒\033[38;5;94;48;5;173m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▓\033[38;5;221;48;5;137m▓\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;101m▒\033[38;5;214;48;5;101m▓\033[38;5;214;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;136;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;165;48;5;230m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;180m░\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m░\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;214;48;5;136m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;136m▒\033[38;5;214;48;5;136m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;222m░\033[38;5;136;48;5;186m░\033[38;5;136;48;5;223m░\033[38;5;136;48;5;222m░\033[38;5;136;48;5;223m░\033[38;5;136;48;5;223m░\033[38;5;178;48;5;223m░\033[38;5;116;48;5;251m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;42;48;5;59m▓\033[38;5;216;48;5;180m░\033[38;5;179;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;179;48;5;136m░\033[38;5;179;48;5;136m░\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;172m▒\033[38;5;179;48;5;172m▒\033[38;5;214;48;5;172m▒\033[38;5;214;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;136m▒\033[38;5;214;48;5;173m▒\033[38;5;179;48;5;172m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;238m▒\033[38;5;221;48;5;237m▒\033[38;5;221;48;5;237m▒\033[38;5;221;48;5;237m▒\033[38;5;221;48;5;237m▒\033[38;5;221;48;5;239m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;136;48;5;223m░\033[38;5;136;48;5;186m░\033[38;5;221;48;5;222m░\033[38;5;136;48;5;223m░\033[38;5;73;48;5;244m▒\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[38;5;131;48;5;236m▒\033[38;5;116;48;5;241m▒\033[38;5;167;48;5;236m░\033[38;5;80;48;5;232m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;80;48;5;234m▒\033[38;5;80;48;5;59m▒\033[38;5;95;48;5;239m▓\033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;7m▒\033[38;5;80;48;5;239m▒\033[38;5;80;48;5;232m▒\033[38;5;209;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;52;48;5;16m \033[38;5;52;48;5;16m \033[38;5;216;48;5;232m \033[38;5;222;48;5;234m \033[38;5;214;48;5;94m░\033[38;5;179;48;5;136m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;173m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;137m▓\033[38;5;136;48;5;240m▒\033[38;5;221;48;5;236m▒\033[38;5;221;48;5;233m░\033[38;5;172;48;5;232m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;52;48;5;16m \033[38;5;136;48;5;232m \033[38;5;221;48;5;235m▒\033[38;5;136;48;5;238m▒\033[38;5;221;48;5;101m▒\033[38;5;221;48;5;101m▒\033[38;5;221;48;5;233m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;136;48;5;234m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;223m░\033[38;5;221;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;51;48;5;230m░\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[0m \033[38;5;138;48;5;238m▓\033[38;5;80;48;5;245m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;131;48;5;238m▒\033[38;5;66;48;5;102m▓\033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;116;48;5;59m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;58m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;143m▓\033[38;5;136;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;236;48;5;236m▓\033[38;5;241;48;5;240m▓\033[38;5;241;48;5;59m▓\033[38;5;235;48;5;234m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;221;48;5;235m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;136;48;5;222m░\033[38;5;221;48;5;186m░\033[38;5;51;48;5;223m░\033[38;5;95;48;5;59m▓\033[0m \033[0m \033[0m \033[0m \033[38;5;95;48;5;240m▓\033[38;5;80;48;5;245m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;234;48;5;234m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;73;48;5;235m▓\033[38;5;66;48;5;243m▓\033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;246m▓\033[38;5;116;48;5;237m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;248;48;5;248m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;232;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;222;48;5;232m \033[38;5;94;48;5;235m▒\033[38;5;94;48;5;58m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;95m▒\033[38;5;136;48;5;237m▒\033[38;5;136;48;5;233m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;221;48;5;232m \033[38;5;136;48;5;236m▒\033[38;5;221;48;5;239m▓\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;144m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;239;48;5;239m▓\033[38;5;247;48;5;246m▓\033[38;5;253;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;249;48;5;249m▓\033[38;5;242;48;5;241m▓\033[38;5;233;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;221;48;5;236m▒\033[38;5;136;48;5;240m▓\033[38;5;221;48;5;236m▒\033[38;5;222;48;5;232m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;221;48;5;232m \033[38;5;94;48;5;236m▒\033[38;5;94;48;5;95m▒\033[38;5;221;48;5;238m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;236m▒\033[38;5;94;48;5;237m▒\033[38;5;214;48;5;232m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;221;48;5;233m▒\033[38;5;221;48;5;237m▒\033[38;5;94;48;5;234m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;88;48;5;238m░\033[38;5;66;48;5;236m▓\033[38;5;242;48;5;242m▓\033[0m \033[0m \033[38;5;95;48;5;240m▓\033[38;5;80;48;5;246m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;249;48;5;249m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;252;48;5;252m▓\033[38;5;233;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;80;48;5;236m░\033[38;5;66;48;5;244m▓\033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;246m▓\033[38;5;73;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;239;48;5;239m▓\033[38;5;246;48;5;246m▓\033[38;5;246;48;5;246m▓\033[38;5;246;48;5;246m▓\033[38;5;246;48;5;246m▓\033[38;5;249;48;5;249m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;7;48;5;7m▓\033[38;5;246;48;5;246m▓\033[38;5;246;48;5;246m▓\033[38;5;246;48;5;246m▓\033[38;5;246;48;5;246m▓\033[38;5;241;48;5;241m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;52;48;5;16m \033[38;5;221;48;5;237m▒\033[38;5;215;48;5;232m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;178;48;5;235m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;178;48;5;101m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;240;48;5;240m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;244;48;5;244m▓\033[38;5;239;48;5;239m▓\033[38;5;239;48;5;239m▓\033[38;5;244;48;5;244m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;243;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;167;48;5;240m░\033[0m \033[0m \033[0m \033[38;5;235;48;5;235m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;246;48;5;246m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;232;48;5;232m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;243;48;5;237m▓\033[38;5;66;48;5;244m▓\033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;109;48;5;243m▓\033[38;5;80;48;5;234m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;237;48;5;237m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;233;48;5;233m▓\033[38;5;7;48;5;250m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;235;48;5;235m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;232;48;5;232m▓\033[38;5;102;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;239;48;5;239m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;221;48;5;95m▓\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;178;48;5;239m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;248;48;5;248m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;237;48;5;237m▓\033[38;5;242;48;5;241m▓\033[38;5;236;48;5;236m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;250;48;5;249m▓\033[38;5;234;48;5;234m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;236;48;5;236m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;80;48;5;254m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;232;48;5;232m▓\033[38;5;250;48;5;250m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;243;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;239;48;5;239m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;167;48;5;240m░\033[0m \033[0m \033[0m \033[38;5;138;48;5;234m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;242;48;5;242m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;249;48;5;249m▓\033[38;5;232;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;95;48;5;238m▓\033[38;5;66;48;5;102m▓\033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;245m▓\033[38;5;66;48;5;241m▓\033[38;5;66;48;5;238m▓\033[38;5;73;48;5;241m▒\033[38;5;116;48;5;233m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;236;48;5;236m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;249;48;5;249m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;241;48;5;59m▓\033[38;5;234;48;5;234m▓\033[38;5;233;48;5;233m▓\033[38;5;240;48;5;240m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;249;48;5;249m▓\033[38;5;232;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;243;48;5;243m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;234;48;5;234m▓\033[38;5;233;48;5;233m▓\033[38;5;237;48;5;237m▓\033[38;5;250;48;5;250m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;233;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;136;48;5;232m░\033[38;5;221;48;5;101m▓\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;137m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;240;48;5;240m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;249;48;5;249m▓\033[38;5;243;48;5;243m▓\033[38;5;239;48;5;238m▓\033[38;5;234;48;5;234m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;247;48;5;247m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;240;48;5;240m▓\033[38;5;233;48;5;233m▓\033[38;5;233;48;5;233m▓\033[38;5;241;48;5;59m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;7;48;5;7m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;247;48;5;247m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;239;48;5;239m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;239;48;5;239m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;253;48;5;253m▓\033[38;5;232;48;5;232m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;249;48;5;249m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;241;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;116;48;5;250m▒\033[0m \033[0m \033[0m \033[38;5;95;48;5;235m▓\033[38;5;37;48;5;232m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;238;48;5;238m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;247m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;80;48;5;59m░\033[38;5;66;48;5;245m▓\033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;241m▓\033[38;5;80;48;5;236m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;236;48;5;236m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;246;48;5;246m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;237;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;232;48;5;233m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;242;48;5;242m▓\033[38;5;16;48;5;16m▓\033[38;5;237;48;5;237m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;251;48;5;251m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;252;48;5;252m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;221;48;5;237m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;239m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;237;48;5;236m▓\033[38;5;247;48;5;247m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;248;48;5;247m▓\033[38;5;234;48;5;234m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;242;48;5;241m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;236;48;5;236m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;237;48;5;237m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;243;48;5;242m▓\033[38;5;16;48;5;16m▓\033[38;5;239;48;5;239m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;248;48;5;247m▓\033[38;5;231;48;5;231m▓\033[38;5;7;48;5;7m▓\033[38;5;239;48;5;238m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;236;48;5;236m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;253;48;5;253m▓\033[38;5;232;48;5;232m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;95;48;5;239m▓\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[0m \033[38;5;95;48;5;236m▓\033[38;5;235;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;246;48;5;246m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;80;48;5;244m▒\033[38;5;66;48;5;247m▓\033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;241m▓\033[38;5;116;48;5;236m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;236;48;5;236m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;248m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;233;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;241;48;5;59m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;248m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;221;48;5;235m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;235m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;232;48;5;233m▓\033[38;5;239;48;5;239m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;235;48;5;235m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;248m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;252;48;5;252m▓\033[38;5;233;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;233;48;5;233m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;247;48;5;247m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;248m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;239;48;5;239m▓\033[38;5;237;48;5;237m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;239;48;5;239m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;248m▓\033[38;5;231;48;5;231m▓\033[38;5;253;48;5;188m▓\033[38;5;236;48;5;236m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;242;48;5;242m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;233;48;5;233m▓\033[38;5;116;48;5;7m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[38;5;238;48;5;238m▓\033[38;5;116;48;5;234m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;233;48;5;233m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;73;48;5;239m▓\033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;241m▓\033[38;5;80;48;5;236m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;237;48;5;237m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;244;48;5;244m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;239;48;5;239m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;237;48;5;237m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;241;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;235;48;5;235m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;235;48;5;235m▓\033[38;5;253;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;249;48;5;249m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;221;48;5;238m▒\033[38;5;221;48;5;95m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;245;48;5;245m▓\033[38;5;249;48;5;249m▓\033[38;5;251;48;5;251m▓\033[38;5;236;48;5;236m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;233;48;5;233m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;238;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;102;48;5;102m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;239;48;5;239m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;237;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;239;48;5;239m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;239m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;237;48;5;237m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;7;48;5;7m▓\033[38;5;252;48;5;252m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;232;48;5;232m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;7;48;5;7m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;80;48;5;102m▒\033[38;5;174;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[38;5;238;48;5;238m▓\033[38;5;80;48;5;234m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;116;48;5;242m▒\033[38;5;174;48;5;235m▒\033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;241m▓\033[38;5;116;48;5;236m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;237;48;5;237m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;245;48;5;245m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;247;48;5;247m▓\033[38;5;241;48;5;59m▓\033[38;5;241;48;5;59m▓\033[38;5;248;48;5;247m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;80;48;5;244m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;238;48;5;238m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;249;48;5;249m▓\033[38;5;242;48;5;241m▓\033[38;5;240;48;5;240m▓\033[38;5;102;48;5;102m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;145;48;5;145m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;136;48;5;234m▒\033[38;5;221;48;5;137m▓\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;232m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;232;48;5;16m▓\033[38;5;247;48;5;247m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;249;48;5;145m▓\033[38;5;246;48;5;246m▓\033[38;5;246;48;5;246m▓\033[38;5;247;48;5;247m▓\033[38;5;251;48;5;251m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;249;48;5;249m▓\033[38;5;232;48;5;232m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;241;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;242;48;5;242m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;246;48;5;246m▓\033[38;5;240;48;5;240m▓\033[38;5;241;48;5;59m▓\033[38;5;248;48;5;248m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;167;48;5;242m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;238;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;246;48;5;246m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;237;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;116;48;5;234m▒\033[38;5;66;48;5;239m▓\033[0m \033[0m \033[0m \033[0m \033[38;5;138;48;5;239m▓\033[38;5;80;48;5;244m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;244;48;5;244m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;232;48;5;232m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;238;48;5;235m▓\033[38;5;66;48;5;242m▓\033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;241m▓\033[38;5;80;48;5;236m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;237;48;5;237m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;243;48;5;242m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;80;48;5;250m░\033[38;5;203;48;5;240m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;238;48;5;238m▓\033[38;5;7;48;5;250m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;253;48;5;253m▓\033[38;5;244;48;5;244m▓\033[38;5;232;48;5;232m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;232m░\033[38;5;118;48;5;137m░\033[38;5;70;48;5;180m▒\033[38;5;35;48;5;180m▒\033[38;5;49;48;5;143m░\033[38;5;220;48;5;233m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;237;48;5;237m▓\033[38;5;249;48;5;249m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;251;48;5;251m▓\033[38;5;242;48;5;241m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;246;48;5;246m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;242;48;5;241m▓\033[38;5;252;48;5;252m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;80;48;5;231m▒\033[38;5;80;48;5;254m░\033[38;5;80;48;5;145m▒\033[38;5;80;48;5;239m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;239;48;5;239m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;109;48;5;250m▓\033[38;5;235;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;236;48;5;236m▓\033[38;5;231;48;5;231m▓\033[38;5;51;48;5;231m \033[38;5;51;48;5;231m \033[38;5;80;48;5;248m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;80;48;5;240m░\033[38;5;95;48;5;239m▓\033[0m \033[0m \033[0m \033[0m \033[38;5;138;48;5;239m▓\033[38;5;80;48;5;242m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;252;48;5;251m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;234;48;5;234m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;80;48;5;234m░\033[38;5;66;48;5;242m▓\033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;244m▓\033[38;5;203;48;5;240m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;244;48;5;237m▓\033[38;5;80;48;5;245m▒\033[38;5;116;48;5;236m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;174;48;5;238m▒\033[38;5;73;48;5;240m▓\033[38;5;247;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;44;48;5;232m░\033[38;5;80;48;5;243m▒\033[38;5;243;48;5;242m▓\033[0m \033[0m \033[0m \033[0m \033[38;5;109;48;5;145m▓\033[38;5;73;48;5;240m▓\033[38;5;43;48;5;235m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;174;48;5;236m▒\033[38;5;181;48;5;239m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;109;48;5;233m▓\033[38;5;116;48;5;245m▒\033[38;5;131;48;5;237m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;238;48;5;237m▓\033[38;5;80;48;5;234m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;116;48;5;243m▒\033[38;5;95;48;5;241m▓\033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;236m▒\033[38;5;116;48;5;246m▒\033[38;5;95;48;5;239m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;167;48;5;236m░\033[38;5;116;48;5;246m▒\033[38;5;131;48;5;236m▒\033[0m \033[0m \033[38;5;131;48;5;237m▓\033[38;5;174;48;5;234m▒\033[38;5;80;48;5;244m▒\033[38;5;167;48;5;236m░\033[38;5;232;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;37;48;5;232m░\033[38;5;167;48;5;238m▒\033[38;5;80;48;5;244m▒\033[38;5;73;48;5;247m▓\033[38;5;167;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;241m▓\033[38;5;80;48;5;246m▒\033[38;5;131;48;5;238m▒\033[38;5;52;48;5;233m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;80;48;5;232m░\033[38;5;131;48;5;236m▒\033[38;5;80;48;5;243m▒\033[38;5;66;48;5;238m▓\033[38;5;95;48;5;239m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;131;48;5;236m▓\033[38;5;116;48;5;245m▒\033[38;5;80;48;5;240m░\033[38;5;80;48;5;234m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;116;48;5;233m▒\033[38;5;167;48;5;238m▒\033[38;5;116;48;5;240m▒\033[38;5;174;48;5;233m▒\033[38;5;138;48;5;238m▓\033[38;5;131;48;5;236m▓\033[38;5;80;48;5;240m▒\033[38;5;80;48;5;232m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;109;48;5;233m▓\033[38;5;80;48;5;244m▒\033[38;5;131;48;5;237m▓\033[38;5;1;48;5;232m░\033[38;5;66;48;5;242m▓\033[38;5;80;48;5;244m▒\033[38;5;73;48;5;235m▓\033[38;5;44;48;5;232m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;44;48;5;232m░\033[38;5;244;48;5;237m▓\033[38;5;80;48;5;244m▒\033[38;5;95;48;5;237m▓\033[38;5;95;48;5;240m▓\033[0m \033[38;5;1;48;5;232m░\033[38;5;66;48;5;241m▓\033[38;5;80;48;5;240m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;116;48;5;234m▒\033[38;5;80;48;5;245m▒\033[38;5;116;48;5;250m▒\033[38;5;80;48;5;59m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;116;48;5;233m▒\033[38;5;80;48;5;243m▒\033[38;5;109;48;5;247m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;235m▒\033[38;5;116;48;5;245m▒\033[38;5;37;48;5;232m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;80;48;5;240m░\033[38;5;80;48;5;252m▒\033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;1;48;5;16m░\033[38;5;1;48;5;16m░\033[38;5;1;48;5;16m░\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
                $display("\033[0m");
			end

			if(err3 == 0) begin
			end
			else if(err4 == 0)
				$display("\n\033[1;32mCongratulations! Your critical path is below 4!\033[m\n");
			else if(err5 == 0)
				$display("\n\033[1;32mCongratulations! Your critical path is below 5!\033[m\n");
			else if(err6 == 0)
				$display("\n\033[1;32mCongratulations! Your critical path is below 6!\033[m\n");
			else if(err7 == 0)
				$display("\n\033[1;32mCongratulations! Your critical path is below 7!\033[m\n");
			else if(err10 == 0)
				$display("\n\033[1;32mCongratulations! Your critical path is below 8!\033[m\n");
			else if(err20 == 0)
				$display("\n\033[1;32mCongratulations! Your score is 40!\033[m\n");
			else begin
			   $display("\nThere are %d errors.\n", err20);
			   $display("Your score is %g.\n", 40-err20/25);
			end

		
			$finish;
		end
		if (err20>100)begin
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;88;48;5;232m░\033[38;5;116;48;5;250m▒\033[38;5;62;48;5;101m▒\033[38;5;220;48;5;240m▓\033[38;5;178;48;5;95m▓\033[38;5;69;48;5;101m░\033[38;5;44;48;5;144m░\033[38;5;80;48;5;253m░\033[38;5;87;48;5;230m░\033[38;5;87;48;5;230m░\033[38;5;87;48;5;230m░\033[38;5;131;48;5;236m▒\033[38;5;131;48;5;236m▒\033[38;5;131;48;5;236m▒\033[38;5;131;48;5;236m▒\033[38;5;131;48;5;236m▒\033[38;5;88;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;239m▓\033[38;5;52;48;5;101m░\033[38;5;221;48;5;94m▒\033[38;5;94;48;5;94m▒\033[38;5;214;48;5;94m▒\033[38;5;179;48;5;94m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;101m▒\033[38;5;172;48;5;101m▓\033[38;5;172;48;5;101m▓\033[38;5;172;48;5;101m▓\033[38;5;130;48;5;101m▓\033[38;5;172;48;5;137m▓\033[38;5;130;48;5;137m▓\033[38;5;172;48;5;137m▓\033[38;5;32;48;5;137m░\033[38;5;26;48;5;137m░\033[38;5;148;48;5;137m▒\033[38;5;209;48;5;144m░\033[38;5;50;48;5;144m░\033[38;5;50;48;5;187m░\033[38;5;50;48;5;187m░\033[38;5;116;48;5;181m▒\033[38;5;35;48;5;242m▓\033[38;5;47;48;5;243m▓\033[38;5;166;48;5;242m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m░\033[38;5;39;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;131m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;94m▒\033[38;5;208;48;5;240m▒\033[38;5;36;48;5;101m░\033[38;5;86;48;5;246m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;224m░\033[38;5;50;48;5;180m░\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;131m▒\033[38;5;130;48;5;130m▒\033[38;5;208;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;208;48;5;58m░\033[38;5;166;48;5;52m \033[38;5;166;48;5;52m \033[38;5;130;48;5;58m \033[38;5;130;48;5;58m░\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;95m▒\033[38;5;130;48;5;95m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;95m▒\033[38;5;172;48;5;58m▒\033[38;5;130;48;5;236m▒\033[38;5;50;48;5;101m░\033[38;5;50;48;5;245m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;238m▓\033[38;5;50;48;5;187m░\033[38;5;179;48;5;143m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;58m░\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;58m \033[38;5;172;48;5;235m \033[38;5;172;48;5;58m▒\033[38;5;50;48;5;101m░\033[38;5;47;48;5;241m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;236m▒\033[38;5;80;48;5;181m░\033[38;5;179;48;5;144m▓\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;95m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;52m \033[38;5;215;48;5;52m \033[38;5;208;48;5;58m░\033[38;5;180;48;5;239m▒\033[38;5;43;48;5;138m▒\033[38;5;49;48;5;245m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m▒\033[38;5;220;48;5;137m▓\033[38;5;172;48;5;144m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;94m░\033[38;5;172;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;208;48;5;130m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;137;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;52m \033[38;5;166;48;5;52m \033[38;5;215;48;5;52m \033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m▒\033[38;5;57;48;5;95m▓\033[38;5;50;48;5;181m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;245m▓\033[38;5;50;48;5;101m▓\033[38;5;220;48;5;59m▓\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;173m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;131m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;95m▒\033[38;5;215;48;5;58m░\033[38;5;202;48;5;52m \033[38;5;216;48;5;52m \033[38;5;166;48;5;52m \033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m▒\033[38;5;166;48;5;58m▒\033[38;5;69;48;5;95m▒\033[38;5;50;48;5;181m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;116;48;5;248m▒\033[38;5;190;48;5;234m▒\033[38;5;58;48;5;234m \033[38;5;172;48;5;95m▒\033[38;5;130;48;5;173m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;130m░\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;95m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;130m▒\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;52m \033[38;5;216;48;5;52m \033[38;5;216;48;5;52m \033[38;5;166;48;5;52m \033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;95m▒\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;246m▒\033[38;5;190;48;5;237m▓\033[38;5;136;48;5;238m▓\033[38;5;137;48;5;95m▒\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;130m▒\033[38;5;172;48;5;136m░\033[38;5;172;48;5;136m░\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;58m▒\033[38;5;76;48;5;238m▓\033[38;5;74;48;5;237m▓\033[38;5;110;48;5;233m▒\033[38;5;137;48;5;232m▓\033[38;5;202;48;5;232m \033[38;5;209;48;5;232m \033[38;5;52;48;5;233m \033[38;5;202;48;5;52m \033[38;5;208;48;5;94m▒\033[38;5;130;48;5;131m▒\033[38;5;130;48;5;137m▒\033[38;5;180;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;130m░\033[38;5;166;48;5;130m░\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;1m░\033[38;5;202;48;5;52m \033[38;5;202;48;5;52m \033[38;5;216;48;5;52m \033[38;5;202;48;5;52m \033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;172;48;5;58m▒\033[38;5;21;48;5;95m░\033[38;5;73;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;101m░\033[38;5;179;48;5;240m▒\033[38;5;179;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;208;48;5;58m░\033[38;5;173;48;5;58m▒\033[38;5;209;48;5;52m▒\033[38;5;204;48;5;239m▓\033[38;5;60;48;5;60m▓\033[38;5;68;48;5;67m▓\033[38;5;26;48;5;66m▓\033[38;5;26;48;5;241m▓\033[38;5;209;48;5;59m▓\033[38;5;166;48;5;95m▓\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;172;48;5;180m░\033[38;5;130;48;5;180m░\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;208;48;5;130m░\033[38;5;180;48;5;130m░\033[38;5;180;48;5;130m░\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;27;48;5;101m▒\033[38;5;80;48;5;253m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;50;48;5;181m▒\033[38;5;121;48;5;240m░\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;208;48;5;94m░\033[38;5;172;48;5;101m▒\033[38;5;220;48;5;101m▓\033[38;5;74;48;5;245m▓\033[38;5;208;48;5;248m▓\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;94;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;180;48;5;130m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;179;48;5;239m▒\033[38;5;176;48;5;101m▒\033[38;5;137;48;5;59m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;16m░\033[38;5;50;48;5;250m▒\033[38;5;94;48;5;101m░\033[38;5;172;48;5;238m▓\033[38;5;172;48;5;236m▒\033[38;5;172;48;5;235m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;131m▒\033[38;5;172;48;5;137m▒\033[38;5;220;48;5;144m▓\033[38;5;25;48;5;246m▓\033[38;5;45;48;5;246m▓\033[38;5;144;48;5;144m▓\033[38;5;220;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;187m▒\033[38;5;214;48;5;187m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;208;48;5;130m▒\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;172;48;5;58m▒\033[38;5;179;48;5;238m▒\033[38;5;21;48;5;59m░\033[38;5;50;48;5;138m▒\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;138;48;5;238m▓\033[38;5;80;48;5;102m░\033[38;5;220;48;5;238m▓\033[38;5;220;48;5;235m▒\033[38;5;220;48;5;235m▒\033[38;5;178;48;5;234m░\033[38;5;214;48;5;235m░\033[38;5;179;48;5;58m░\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;101m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;94;48;5;144m▓\033[38;5;39;48;5;109m▓\033[38;5;25;48;5;67m▓\033[38;5;35;48;5;248m▓\033[38;5;112;48;5;151m▓\033[38;5;190;48;5;187m▓\033[38;5;144;48;5;187m▓\033[38;5;178;48;5;187m▓\033[38;5;178;48;5;187m▓\033[38;5;214;48;5;188m▓\033[38;5;179;48;5;188m▒\033[38;5;172;48;5;187m▒\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;95m▓\033[38;5;50;48;5;181m░\033[38;5;86;48;5;246m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;145m▓\033[38;5;216;48;5;239m░\033[38;5;58;48;5;232m \033[38;5;58;48;5;232m \033[38;5;58;48;5;233m \033[38;5;58;48;5;233m \033[38;5;220;48;5;233m \033[38;5;136;48;5;235m░\033[38;5;221;48;5;58m▒\033[38;5;179;48;5;95m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;101m▒\033[38;5;214;48;5;101m▒\033[38;5;94;48;5;137m▒\033[38;5;112;48;5;244m▓\033[38;5;39;48;5;60m▓\033[38;5;35;48;5;245m▓\033[38;5;190;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;172;48;5;181m▓\033[38;5;179;48;5;187m▓\033[38;5;130;48;5;187m▒\033[38;5;130;48;5;187m▒\033[38;5;130;48;5;187m▒\033[38;5;172;48;5;187m▒\033[38;5;172;48;5;187m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;208;48;5;58m▒\033[38;5;172;48;5;95m▓\033[38;5;80;48;5;181m▒\033[38;5;43;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;131;48;5;240m▓\033[38;5;143;48;5;232m▒\033[38;5;58;48;5;232m \033[38;5;190;48;5;232m \033[38;5;220;48;5;232m \033[38;5;136;48;5;232m \033[38;5;222;48;5;232m \033[38;5;172;48;5;233m \033[38;5;221;48;5;235m░\033[38;5;94;48;5;240m▒\033[38;5;214;48;5;101m▓\033[38;5;172;48;5;101m▒\033[38;5;172;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;214;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;221;48;5;94m▒\033[38;5;220;48;5;58m▒\033[38;5;143;48;5;237m▒\033[38;5;178;48;5;239m▓\033[38;5;221;48;5;95m▓\033[38;5;179;48;5;137m▓\033[38;5;214;48;5;144m▓\033[38;5;136;48;5;144m▓\033[38;5;221;48;5;144m▒\033[38;5;221;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;131m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;221;48;5;58m▒\033[38;5;221;48;5;95m▓\033[38;5;50;48;5;144m░\033[38;5;149;48;5;59m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;116;48;5;246m▒\033[38;5;190;48;5;233m▓\033[38;5;155;48;5;16m \033[38;5;58;48;5;232m \033[38;5;220;48;5;232m \033[38;5;136;48;5;232m \033[38;5;214;48;5;232m \033[38;5;136;48;5;234m░\033[38;5;221;48;5;238m▒\033[38;5;94;48;5;95m▓\033[38;5;179;48;5;101m▓\033[38;5;214;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;94m▒\033[38;5;221;48;5;58m▒\033[38;5;178;48;5;58m░\033[38;5;172;48;5;234m \033[38;5;172;48;5;233m \033[38;5;221;48;5;58m░\033[38;5;221;48;5;95m▒\033[38;5;221;48;5;101m▓\033[38;5;94;48;5;143m▓\033[38;5;221;48;5;144m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;143m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;131m▒\033[38;5;180;48;5;130m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;179;48;5;94m▒\033[38;5;214;48;5;94m▒\033[38;5;94;48;5;94m▒\033[38;5;94;48;5;95m▒\033[38;5;50;48;5;144m░\033[38;5;49;48;5;243m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;241;48;5;240m▓\033[38;5;80;48;5;242m▒\033[38;5;143;48;5;235m▓\033[38;5;220;48;5;235m▒\033[38;5;220;48;5;235m▒\033[38;5;220;48;5;235m▒\033[38;5;178;48;5;236m▒\033[38;5;221;48;5;238m▓\033[38;5;94;48;5;59m▓\033[38;5;214;48;5;95m▓\033[38;5;214;48;5;95m▒\033[38;5;94;48;5;58m▒\033[38;5;221;48;5;58m▒\033[38;5;221;48;5;58m▒\033[38;5;221;48;5;58m░\033[38;5;222;48;5;234m \033[38;5;94;48;5;234m \033[38;5;136;48;5;58m░\033[38;5;221;48;5;58m▒\033[38;5;136;48;5;95m▒\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;137m▓\033[38;5;94;48;5;144m▓\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;131m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;214;48;5;94m▒\033[38;5;221;48;5;94m▒\033[38;5;221;48;5;95m▒\033[38;5;80;48;5;181m▒\033[38;5;50;48;5;246m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;109;48;5;248m▓\033[38;5;66;48;5;244m▓\033[38;5;109;48;5;241m▓\033[38;5;116;48;5;243m▒\033[38;5;80;48;5;243m▒\033[38;5;220;48;5;59m▒\033[38;5;136;48;5;238m▒\033[38;5;178;48;5;58m▒\033[38;5;178;48;5;58m▒\033[38;5;178;48;5;58m▒\033[38;5;178;48;5;58m░\033[38;5;136;48;5;58m▒\033[38;5;136;48;5;240m▒\033[38;5;136;48;5;101m▒\033[38;5;221;48;5;101m▓\033[38;5;136;48;5;101m▓\033[38;5;221;48;5;137m▓\033[38;5;136;48;5;143m▓\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;131m▒\033[38;5;180;48;5;130m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;179;48;5;94m▒\033[38;5;94;48;5;94m▒\033[38;5;136;48;5;94m▒\033[38;5;178;48;5;94m▒\033[38;5;33;48;5;101m▒\033[38;5;80;48;5;187m░\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▒\033[38;5;80;48;5;144m▒\033[38;5;220;48;5;101m▓\033[38;5;178;48;5;101m▓\033[38;5;178;48;5;101m▒\033[38;5;136;48;5;95m▒\033[38;5;136;48;5;101m▓\033[38;5;221;48;5;101m▓\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;143m▓\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;216;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;179;48;5;94m▒\033[38;5;214;48;5;95m▒\033[38;5;50;48;5;144m░\033[38;5;131;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m▒\033[38;5;220;48;5;101m▓\033[38;5;178;48;5;101m▓\033[38;5;221;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;214;48;5;137m▓\033[38;5;214;48;5;137m▓\033[38;5;179;48;5;144m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;216;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;215;48;5;94m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;130;48;5;95m▒\033[38;5;55;48;5;138m▒\033[38;5;50;48;5;144m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;252m▒\033[38;5;220;48;5;144m▓\033[38;5;136;48;5;144m▓\033[38;5;214;48;5;144m▓\033[38;5;179;48;5;144m▓\033[38;5;172;48;5;144m▓\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;131m▒\033[38;5;180;48;5;130m▒\033[38;5;180;48;5;130m▒\033[38;5;166;48;5;94m▒\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m▒\033[38;5;130;48;5;95m▒\033[38;5;84;48;5;138m▒\033[38;5;86;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;252m▒\033[38;5;178;48;5;144m▓\033[38;5;214;48;5;144m▓\033[38;5;172;48;5;144m▓\033[38;5;130;48;5;144m▓\033[38;5;130;48;5;144m▓\033[38;5;130;48;5;144m▓\033[38;5;130;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;144m▒\033[38;5;179;48;5;144m▒\033[38;5;221;48;5;144m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;180;48;5;130m▒\033[38;5;180;48;5;130m▒\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;180;48;5;130m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;208;48;5;58m▒\033[38;5;172;48;5;95m▒\033[38;5;226;48;5;144m░\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;252m▒\033[38;5;214;48;5;249m▓\033[38;5;172;48;5;180m▓\033[38;5;172;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▓\033[38;5;130;48;5;180m▓\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;144m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;180;48;5;130m░\033[38;5;180;48;5;130m░\033[38;5;166;48;5;130m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;173;48;5;94m░\033[38;5;202;48;5;94m░\033[38;5;173;48;5;94m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;94m░\033[38;5;202;48;5;94m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;208;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;202;48;5;52m░\033[38;5;166;48;5;58m░\033[38;5;180;48;5;94m░\033[38;5;208;48;5;94m▒\033[38;5;172;48;5;95m▓\033[38;5;80;48;5;144m░\033[38;5;131;48;5;237m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;252m▒\033[38;5;172;48;5;249m▓\033[38;5;172;48;5;95m▓\033[38;5;130;48;5;234m▓\033[38;5;130;48;5;234m▓\033[38;5;130;48;5;234m▓\033[38;5;172;48;5;234m▓\033[38;5;130;48;5;234m▓\033[38;5;130;48;5;234m▓\033[38;5;172;48;5;234m▓\033[38;5;172;48;5;234m▓\033[38;5;130;48;5;234m▓\033[38;5;130;48;5;234m▓\033[38;5;214;48;5;234m▓\033[38;5;94;48;5;234m▒\033[38;5;221;48;5;233m▒\033[38;5;222;48;5;233m░\033[38;5;179;48;5;236m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;58m░\033[38;5;209;48;5;232m \033[38;5;209;48;5;232m \033[38;5;209;48;5;232m \033[38;5;209;48;5;232m \033[38;5;209;48;5;232m \033[38;5;202;48;5;233m \033[38;5;180;48;5;94m░\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;234m░\033[38;5;216;48;5;232m \033[38;5;216;48;5;232m \033[38;5;202;48;5;233m \033[38;5;202;48;5;232m \033[38;5;215;48;5;234m░\033[38;5;180;48;5;58m▒\033[38;5;208;48;5;234m░\033[38;5;202;48;5;232m \033[38;5;216;48;5;232m \033[38;5;209;48;5;232m \033[38;5;216;48;5;232m \033[38;5;130;48;5;234m░\033[38;5;208;48;5;58m░\033[38;5;208;48;5;94m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;202;48;5;52m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m░\033[38;5;180;48;5;94m▒\033[38;5;130;48;5;95m▒\033[38;5;43;48;5;101m░\033[38;5;50;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;116;48;5;246m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;137m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;215;48;5;52m░\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;172;48;5;95m▒\033[38;5;50;48;5;180m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;238;48;5;238m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;172;48;5;236m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;234m \033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;52m░\033[38;5;166;48;5;52m░\033[38;5;166;48;5;52m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;62;48;5;101m▒\033[38;5;50;48;5;144m▓\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;238m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;252;48;5;252m▓\033[38;5;252;48;5;252m▓\033[38;5;252;48;5;252m▓\033[38;5;252;48;5;252m▓\033[38;5;252;48;5;252m▓\033[38;5;252;48;5;252m▓\033[38;5;252;48;5;252m▓\033[38;5;252;48;5;252m▓\033[38;5;240;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;235;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;253;48;5;253m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;52;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;234m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;52m░\033[38;5;202;48;5;52m \033[38;5;202;48;5;52m \033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;58m▒\033[38;5;201;48;5;101m░\033[38;5;29;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;238m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;188;48;5;252m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;240m▓\033[38;5;249;48;5;249m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;234m░\033[38;5;166;48;5;94m▒\033[38;5;202;48;5;58m░\033[38;5;202;48;5;52m░\033[38;5;216;48;5;52m \033[38;5;216;48;5;52m \033[38;5;166;48;5;52m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m▒\033[38;5;50;48;5;144m▒\033[38;5;131;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;238m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;248;48;5;248m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;237;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;235m░\033[38;5;166;48;5;94m░\033[38;5;202;48;5;52m░\033[38;5;216;48;5;52m \033[38;5;216;48;5;52m \033[38;5;166;48;5;52m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;52m░\033[38;5;179;48;5;236m▒\033[38;5;80;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;237m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;234;48;5;234m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;235;48;5;235m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;232;48;5;232m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;238;48;5;238m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;234m \033[38;5;166;48;5;58m░\033[38;5;166;48;5;52m░\033[38;5;202;48;5;52m \033[38;5;202;48;5;52m \033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;208;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;208;48;5;52m \033[38;5;130;48;5;234m░\033[38;5;190;48;5;239m░\033[38;5;109;48;5;248m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;243;48;5;243m▓\033[38;5;73;48;5;237m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;7;48;5;7m▓\033[38;5;7;48;5;7m▓\033[38;5;251;48;5;251m▓\033[38;5;7;48;5;7m▓\033[38;5;7;48;5;7m▓\033[38;5;7;48;5;7m▓\033[38;5;251;48;5;251m▓\033[38;5;7;48;5;7m▓\033[38;5;232;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;252;48;5;252m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;209;48;5;232m \033[38;5;202;48;5;52m \033[38;5;216;48;5;234m \033[38;5;216;48;5;234m \033[38;5;202;48;5;52m \033[38;5;166;48;5;52m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m░\033[38;5;208;48;5;58m░\033[38;5;166;48;5;52m \033[38;5;166;48;5;52m \033[38;5;215;48;5;52m \033[38;5;208;48;5;235m░\033[38;5;130;48;5;234m░\033[38;5;50;48;5;243m▒\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;237m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;249;48;5;249m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;238;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;52;48;5;16m \033[38;5;166;48;5;94m░\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;215;48;5;58m░\033[38;5;215;48;5;52m \033[38;5;166;48;5;52m \033[38;5;166;48;5;52m \033[38;5;166;48;5;52m \033[38;5;166;48;5;52m \033[38;5;215;48;5;52m░\033[38;5;84;48;5;236m▒\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;243;48;5;242m▓\033[38;5;50;48;5;237m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;237m▓\033[38;5;179;48;5;240m▓\033[38;5;172;48;5;236m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;242;48;5;241m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;233;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;239;48;5;239m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;233;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;248;48;5;247m▓\033[38;5;248;48;5;247m▓\033[38;5;248;48;5;247m▓\033[38;5;248;48;5;247m▓\033[38;5;248;48;5;247m▓\033[38;5;248;48;5;247m▓\033[38;5;248;48;5;247m▓\033[38;5;248;48;5;247m▓\033[38;5;243;48;5;242m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;52m░\033[38;5;166;48;5;94m░\033[38;5;180;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;52m \033[38;5;166;48;5;52m \033[38;5;166;48;5;52m \033[38;5;166;48;5;52m \033[38;5;215;48;5;52m \033[38;5;208;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;50;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;244;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;172;48;5;101m▓\033[38;5;179;48;5;144m▓\033[38;5;52;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;238;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;214;48;5;235m▒\033[38;5;94;48;5;233m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;248;48;5;248m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;252;48;5;252m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;7;48;5;7m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;234m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;52m░\033[38;5;166;48;5;52m \033[38;5;215;48;5;52m░\033[38;5;215;48;5;52m░\033[38;5;215;48;5;58m░\033[38;5;208;48;5;58m▒\033[38;5;172;48;5;240m▒\033[38;5;50;48;5;101m░\033[38;5;47;48;5;243m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;73;48;5;245m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;232m \033[38;5;179;48;5;144m▓\033[38;5;179;48;5;144m▒\033[38;5;179;48;5;234m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;238m▓\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;233m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;208;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;45;48;5;240m▒\033[38;5;202;48;5;241m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;253m░\033[38;5;76;48;5;144m░\033[38;5;221;48;5;237m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;232m \033[38;5;136;48;5;101m▓\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;144m▓\033[38;5;179;48;5;234m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;221;48;5;237m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;234m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;52;48;5;16m \033[38;5;215;48;5;233m \033[38;5;52;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;52;48;5;16m \033[38;5;215;48;5;52m░\033[38;5;180;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;45;48;5;238m░\033[38;5;209;48;5;59m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;254m░\033[38;5;162;48;5;144m▒\033[38;5;136;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;136;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m▒\033[38;5;38;48;5;240m▒\033[38;5;202;48;5;241m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;70;48;5;143m░\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;50;48;5;101m▒\033[38;5;174;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;55;48;5;137m▓\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;143m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;180;48;5;58m░\033[38;5;208;48;5;58m▒\033[38;5;208;48;5;237m▒\033[38;5;69;48;5;239m░\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;254m░\033[38;5;76;48;5;137m░\033[38;5;221;48;5;101m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;208;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m \033[38;5;130;48;5;58m░\033[38;5;130;48;5;52m░\033[38;5;130;48;5;236m░\033[38;5;130;48;5;236m▒\033[38;5;209;48;5;240m▒\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;254m░\033[38;5;119;48;5;137m░\033[38;5;221;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;208;48;5;58m░\033[38;5;215;48;5;52m \033[38;5;215;48;5;52m \033[38;5;130;48;5;52m \033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;208;48;5;58m▒\033[38;5;130;48;5;237m▒\033[38;5;82;48;5;238m▒\033[38;5;49;48;5;242m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;254m░\033[38;5;46;48;5;137m░\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;208;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;215;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;215;48;5;52m \033[38;5;215;48;5;52m \033[38;5;215;48;5;52m \033[38;5;130;48;5;52m \033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;130;48;5;58m▒\033[38;5;77;48;5;238m▒\033[38;5;50;48;5;247m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;254m░\033[38;5;46;48;5;137m░\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;143m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;95m▒\033[38;5;214;48;5;94m▒\033[38;5;94;48;5;94m▒\033[38;5;94;48;5;94m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;221;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;101m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;208;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;166;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m░\033[38;5;215;48;5;58m░\033[38;5;215;48;5;52m \033[38;5;215;48;5;52m \033[38;5;166;48;5;234m \033[38;5;215;48;5;52m \033[38;5;208;48;5;52m \033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;130;48;5;58m▒\033[38;5;130;48;5;58m▒\033[38;5;130;48;5;58m▒\033[38;5;70;48;5;95m░\033[38;5;50;48;5;181m▒\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;253m░\033[38;5;32;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;94m▒\033[38;5;214;48;5;58m░\033[38;5;214;48;5;58m \033[38;5;214;48;5;58m \033[38;5;94;48;5;58m▒\033[38;5;94;48;5;95m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;214;48;5;94m▒\033[38;5;179;48;5;136m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;208;48;5;130m▒\033[38;5;180;48;5;94m░\033[38;5;180;48;5;94m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;215;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;52m \033[38;5;215;48;5;234m \033[38;5;166;48;5;234m \033[38;5;166;48;5;234m \033[38;5;215;48;5;52m \033[38;5;130;48;5;52m \033[38;5;130;48;5;52m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;208;48;5;58m░\033[38;5;104;48;5;95m▒\033[38;5;42;48;5;101m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;138;48;5;239m▓\033[38;5;109;48;5;247m▓\033[38;5;80;48;5;187m░\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;95m▒\033[38;5;136;48;5;58m▒\033[38;5;221;48;5;58m \033[38;5;214;48;5;235m \033[38;5;222;48;5;235m \033[38;5;214;48;5;58m \033[38;5;94;48;5;58m░\033[38;5;214;48;5;94m▒\033[38;5;214;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;214;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;180;48;5;130m▒\033[38;5;180;48;5;130m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;130;48;5;58m░\033[38;5;172;48;5;52m \033[38;5;215;48;5;234m \033[38;5;166;48;5;233m \033[38;5;166;48;5;234m \033[38;5;215;48;5;234m \033[38;5;130;48;5;52m \033[38;5;172;48;5;52m░\033[38;5;172;48;5;58m░\033[38;5;222;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;236m▒\033[38;5;36;48;5;95m▒\033[38;5;174;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;109;48;5;247m▓\033[38;5;109;48;5;246m▓\033[38;5;80;48;5;188m░\033[38;5;208;48;5;250m▒\033[38;5;101;48;5;144m▓\033[38;5;144;48;5;143m▓\033[38;5;220;48;5;143m▓\033[38;5;221;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;178;48;5;101m▒\033[38;5;178;48;5;58m▒\033[38;5;178;48;5;58m▒\033[38;5;178;48;5;58m░\033[38;5;178;48;5;58m░\033[38;5;221;48;5;58m░\033[38;5;94;48;5;58m░\033[38;5;214;48;5;58m░\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;95m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;173m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;208;48;5;130m▒\033[38;5;180;48;5;130m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;52m \033[38;5;166;48;5;234m \033[38;5;166;48;5;233m \033[38;5;130;48;5;234m \033[38;5;172;48;5;234m \033[38;5;222;48;5;235m \033[38;5;222;48;5;235m \033[38;5;214;48;5;235m \033[38;5;214;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;222;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;56;48;5;238m░\033[38;5;72;48;5;59m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;254m░\033[38;5;80;48;5;187m░\033[38;5;44;48;5;187m░\033[38;5;29;48;5;144m░\033[38;5;144;48;5;101m▓\033[38;5;144;48;5;101m▓\033[38;5;144;48;5;101m▓\033[38;5;143;48;5;101m▓\033[38;5;143;48;5;101m▓\033[38;5;143;48;5;101m▓\033[38;5;220;48;5;101m▒\033[38;5;220;48;5;101m▒\033[38;5;136;48;5;137m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;178;48;5;137m▓\033[38;5;220;48;5;94m▒\033[38;5;220;48;5;58m▒\033[38;5;178;48;5;58m░\033[38;5;178;48;5;58m░\033[38;5;136;48;5;58m░\033[38;5;221;48;5;235m░\033[38;5;222;48;5;234m \033[38;5;222;48;5;235m░\033[38;5;179;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;179;48;5;95m▒\033[38;5;94;48;5;101m▒\033[38;5;214;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;173m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;130m▒\033[38;5;208;48;5;130m▒\033[38;5;208;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;130;48;5;52m \033[38;5;166;48;5;234m \033[38;5;166;48;5;234m \033[38;5;130;48;5;234m \033[38;5;172;48;5;234m \033[38;5;222;48;5;235m \033[38;5;214;48;5;235m \033[38;5;214;48;5;235m \033[38;5;222;48;5;235m░\033[38;5;222;48;5;58m░\033[38;5;222;48;5;58m░\033[38;5;214;48;5;58m░\033[38;5;222;48;5;58m░\033[38;5;214;48;5;58m░\033[38;5;222;48;5;58m░\033[38;5;222;48;5;58m░\033[38;5;77;48;5;58m░\033[38;5;86;48;5;101m▒\033[38;5;167;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;236m▒\033[38;5;87;48;5;254m░\033[38;5;44;48;5;187m░\033[38;5;77;48;5;144m░\033[38;5;220;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;144;48;5;144m▓\033[38;5;220;48;5;143m▓\033[38;5;220;48;5;137m▓\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;101m▒\033[38;5;143;48;5;95m▒\033[38;5;220;48;5;240m▒\033[38;5;220;48;5;58m▒\033[38;5;220;48;5;58m▒\033[38;5;220;48;5;58m▒\033[38;5;220;48;5;94m▒\033[38;5;221;48;5;101m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;178;48;5;143m▒\033[38;5;178;48;5;143m▒\033[38;5;220;48;5;101m▒\033[38;5;178;48;5;94m▒\033[38;5;178;48;5;58m░\033[38;5;136;48;5;58m░\033[38;5;136;48;5;58m \033[38;5;222;48;5;234m \033[38;5;172;48;5;234m \033[38;5;94;48;5;235m \033[38;5;214;48;5;58m▒\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;101m▓\033[38;5;221;48;5;101m▓\033[38;5;94;48;5;101m▓\033[38;5;214;48;5;137m▓\033[38;5;221;48;5;137m▓\033[38;5;221;48;5;101m▓\033[38;5;221;48;5;101m▓\033[38;5;94;48;5;101m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;131m▒\033[38;5;208;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;52m░\033[38;5;166;48;5;234m \033[38;5;215;48;5;234m \033[38;5;130;48;5;234m \033[38;5;172;48;5;234m \033[38;5;172;48;5;235m \033[38;5;222;48;5;235m \033[38;5;214;48;5;235m░\033[38;5;222;48;5;235m░\033[38;5;222;48;5;236m░\033[38;5;222;48;5;235m░\033[38;5;222;48;5;235m \033[38;5;94;48;5;235m \033[38;5;221;48;5;235m░\033[38;5;77;48;5;235m░\033[38;5;50;48;5;95m▒\033[38;5;209;48;5;237m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;253m░\033[38;5;178;48;5;144m▓\033[38;5;220;48;5;144m▓\033[38;5;144;48;5;143m▓\033[38;5;144;48;5;143m▓\033[38;5;144;48;5;137m▓\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;95m▓\033[38;5;178;48;5;95m▓\033[38;5;178;48;5;95m▓\033[38;5;220;48;5;240m▓\033[38;5;178;48;5;240m▓\033[38;5;84;48;5;240m░\033[38;5;80;48;5;101m░\033[38;5;50;48;5;144m▒\033[38;5;50;48;5;180m▒\033[38;5;50;48;5;143m░\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;137m▒\033[38;5;178;48;5;101m▒\033[38;5;220;48;5;58m▒\033[38;5;178;48;5;58m▒\033[38;5;136;48;5;58m░\033[38;5;136;48;5;58m░\033[38;5;221;48;5;58m▒\033[38;5;221;48;5;95m▒\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;101m▓\033[38;5;136;48;5;101m▓\033[38;5;214;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;136;48;5;137m▓\033[38;5;221;48;5;137m▓\033[38;5;221;48;5;137m▓\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;130;48;5;131m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;52m░\033[38;5;166;48;5;234m \033[38;5;215;48;5;234m \033[38;5;130;48;5;234m \033[38;5;172;48;5;234m \033[38;5;172;48;5;234m \033[38;5;172;48;5;235m \033[38;5;222;48;5;235m \033[38;5;222;48;5;235m░\033[38;5;214;48;5;235m░\033[38;5;222;48;5;235m░\033[38;5;130;48;5;233m \033[38;5;161;48;5;234m▓\033[38;5;43;48;5;101m▓\033[38;5;131;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;246m▒\033[38;5;220;48;5;235m▒\033[38;5;144;48;5;240m▓\033[38;5;144;48;5;101m▓\033[38;5;143;48;5;240m▒\033[38;5;185;48;5;235m░\033[38;5;185;48;5;236m▒\033[38;5;143;48;5;240m▓\033[38;5;130;48;5;241m░\033[38;5;80;48;5;101m░\033[38;5;116;48;5;144m▒\033[38;5;66;48;5;102m▓\033[38;5;174;48;5;234m▒\033[38;5;174;48;5;235m▒\033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;43;48;5;180m░\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;136;48;5;101m▒\033[38;5;178;48;5;58m▒\033[38;5;220;48;5;58m▒\033[38;5;178;48;5;58m▒\033[38;5;136;48;5;58m▒\033[38;5;136;48;5;95m▒\033[38;5;136;48;5;101m▒\033[38;5;221;48;5;101m▓\033[38;5;94;48;5;137m▓\033[38;5;179;48;5;137m▓\033[38;5;179;48;5;137m▓\033[38;5;179;48;5;137m▓\033[38;5;179;48;5;137m▓\033[38;5;179;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;214;48;5;137m▓\033[38;5;94;48;5;143m▓\033[38;5;136;48;5;143m▓\033[38;5;136;48;5;143m▓\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;58m░\033[38;5;215;48;5;234m \033[38;5;208;48;5;234m \033[38;5;130;48;5;234m \033[38;5;130;48;5;234m \033[38;5;172;48;5;234m \033[38;5;222;48;5;234m \033[38;5;222;48;5;234m \033[38;5;222;48;5;234m \033[38;5;179;48;5;235m░\033[38;5;218;48;5;238m░\033[38;5;42;48;5;242m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;138;48;5;239m▓\033[38;5;73;48;5;249m▒\033[38;5;73;48;5;246m▓\033[38;5;116;48;5;250m▒\033[38;5;73;48;5;246m▓\033[38;5;109;48;5;243m▓\033[38;5;109;48;5;244m▓\033[38;5;73;48;5;250m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m▒\033[38;5;83;48;5;137m░\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;101m▒\033[38;5;221;48;5;94m▒\033[38;5;136;48;5;58m▒\033[38;5;136;48;5;58m░\033[38;5;178;48;5;58m▒\033[38;5;178;48;5;58m▒\033[38;5;178;48;5;94m▒\033[38;5;136;48;5;101m▒\033[38;5;136;48;5;101m▓\033[38;5;221;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;144m▓\033[38;5;172;48;5;144m▓\033[38;5;172;48;5;144m▓\033[38;5;179;48;5;144m▓\033[38;5;172;48;5;144m▓\033[38;5;172;48;5;144m▓\033[38;5;172;48;5;144m▓\033[38;5;214;48;5;144m▓\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;235m \033[38;5;215;48;5;234m \033[38;5;215;48;5;233m \033[38;5;130;48;5;233m \033[38;5;172;48;5;234m \033[38;5;172;48;5;233m \033[38;5;172;48;5;235m▒\033[38;5;103;48;5;236m▓\033[38;5;36;48;5;95m▒\033[38;5;50;48;5;145m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;86;48;5;95m▓\033[38;5;76;48;5;101m░\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;100m▒\033[38;5;221;48;5;94m▒\033[38;5;136;48;5;58m░\033[38;5;178;48;5;58m░\033[38;5;220;48;5;58m░\033[38;5;178;48;5;94m▒\033[38;5;178;48;5;101m▒\033[38;5;136;48;5;137m▓\033[38;5;136;48;5;143m▓\033[38;5;221;48;5;143m▓\033[38;5;94;48;5;144m▓\033[38;5;94;48;5;144m▓\033[38;5;214;48;5;144m▓\033[38;5;179;48;5;144m▓\033[38;5;179;48;5;144m▓\033[38;5;179;48;5;144m▓\033[38;5;179;48;5;144m▒\033[38;5;172;48;5;144m▒\033[38;5;172;48;5;144m▓\033[38;5;94;48;5;144m▓\033[38;5;221;48;5;143m▓\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;234m \033[38;5;166;48;5;233m \033[38;5;215;48;5;233m \033[38;5;166;48;5;233m \033[38;5;130;48;5;233m \033[38;5;112;48;5;236m░\033[38;5;43;48;5;59m▓\033[38;5;84;48;5;243m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;235m▒\033[38;5;79;48;5;243m▓\033[38;5;73;48;5;144m▒\033[38;5;80;48;5;144m▒\033[38;5;31;48;5;101m▓\033[38;5;221;48;5;101m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;136;48;5;137m▒\033[38;5;221;48;5;136m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;101m▒\033[38;5;94;48;5;94m▒\033[38;5;221;48;5;58m▒\033[38;5;136;48;5;58m▒\033[38;5;178;48;5;101m▒\033[38;5;136;48;5;137m▓\033[38;5;221;48;5;144m▓\033[38;5;221;48;5;144m▒\033[38;5;94;48;5;144m▓\033[38;5;94;48;5;144m▓\033[38;5;214;48;5;144m▓\033[38;5;94;48;5;144m▓\033[38;5;214;48;5;144m▓\033[38;5;214;48;5;144m▓\033[38;5;179;48;5;144m▓\033[38;5;179;48;5;144m▓\033[38;5;94;48;5;144m▓\033[38;5;94;48;5;144m▓\033[38;5;94;48;5;144m▓\033[38;5;221;48;5;137m▓\033[38;5;136;48;5;137m▓\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;130;48;5;236m░\033[38;5;166;48;5;233m \033[38;5;166;48;5;233m \033[38;5;174;48;5;237m▒\033[38;5;220;48;5;238m▓\033[38;5;174;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;249m▒\033[38;5;116;48;5;144m▒\033[38;5;80;48;5;181m░\033[38;5;153;48;5;144m░\033[38;5;81;48;5;101m░\033[38;5;94;48;5;101m▓\033[38;5;214;48;5;95m▓\033[38;5;179;48;5;95m▒\033[38;5;94;48;5;94m▒\033[38;5;221;48;5;3m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;137m▒\033[38;5;136;48;5;101m▒\033[38;5;50;48;5;137m░\033[38;5;50;48;5;137m▒\033[38;5;50;48;5;101m░\033[38;5;29;48;5;95m▓\033[38;5;32;48;5;101m▒\033[38;5;27;48;5;138m▒\033[38;5;57;48;5;144m░\033[38;5;94;48;5;181m▓\033[38;5;136;48;5;181m▓\033[38;5;94;48;5;181m▓\033[38;5;94;48;5;181m▓\033[38;5;94;48;5;181m▓\033[38;5;179;48;5;180m▓\033[38;5;221;48;5;144m▓\033[38;5;94;48;5;144m▓\033[38;5;221;48;5;144m▓\033[38;5;136;48;5;144m▓\033[38;5;178;48;5;144m▓\033[38;5;136;48;5;137m▓\033[38;5;178;48;5;101m▓\033[38;5;178;48;5;95m▓\033[38;5;221;48;5;58m▒\033[38;5;94;48;5;101m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;208;48;5;58m░\033[38;5;180;48;5;58m▒\033[38;5;180;48;5;237m▒\033[38;5;137;48;5;237m▒\033[38;5;50;48;5;241m▒\033[38;5;50;48;5;248m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;254m░\033[38;5;171;48;5;101m░\033[38;5;119;48;5;101m░\033[38;5;178;48;5;101m▓\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;101m▓\033[38;5;221;48;5;101m▓\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;101m▒\033[38;5;136;48;5;101m▒\033[38;5;136;48;5;101m▒\033[38;5;221;48;5;95m▒\033[38;5;221;48;5;95m▒\033[38;5;136;48;5;101m▒\033[38;5;178;48;5;137m▒\033[38;5;178;48;5;143m▒\033[38;5;178;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;178;48;5;137m▓\033[38;5;50;48;5;144m▒\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;116;48;5;187m▒\033[38;5;73;48;5;144m▒\033[38;5;50;48;5;137m▒\033[38;5;110;48;5;95m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;180;48;5;58m▒\033[38;5;208;48;5;236m▒\033[38;5;43;48;5;240m░\033[38;5;209;48;5;239m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;246m▓\033[38;5;21;48;5;238m░\033[38;5;220;48;5;233m \033[38;5;220;48;5;235m░\033[38;5;136;48;5;58m▒\033[38;5;136;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;101m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;178;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;112;48;5;143m▒\033[38;5;73;48;5;246m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;236m▒\033[38;5;50;48;5;180m░\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;180;48;5;58m▒\033[38;5;43;48;5;95m░\033[38;5;86;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;246m▓\033[38;5;93;48;5;101m░\033[38;5;136;48;5;101m▓\033[38;5;178;48;5;101m▓\033[38;5;178;48;5;137m▓\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;220;48;5;179m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;86;48;5;143m░\033[38;5;80;48;5;186m▒\033[38;5;131;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;236m▒\033[38;5;50;48;5;180m░\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;208;48;5;58m░\033[38;5;38;48;5;239m▓\033[38;5;36;48;5;138m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;7m▒\033[38;5;45;48;5;95m░\033[38;5;136;48;5;101m▓\033[38;5;178;48;5;137m▒\033[38;5;136;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;178;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▓\033[38;5;80;48;5;187m░\033[38;5;131;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;236m▒\033[38;5;50;48;5;187m░\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;215;48;5;58m░\033[38;5;36;48;5;95m░\033[38;5;50;48;5;249m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;187m▒\033[38;5;44;48;5;187m░\033[38;5;220;48;5;137m▓\033[38;5;220;48;5;137m▓\033[38;5;220;48;5;143m▒\033[38;5;178;48;5;143m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;201;48;5;144m░\033[38;5;50;48;5;187m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;230m░\033[38;5;104;48;5;180m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m▒\033[38;5;200;48;5;95m▒\033[38;5;50;48;5;248m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;138;48;5;238m▓\033[38;5;80;48;5;144m▒\033[38;5;84;48;5;101m░\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;137m▓\033[38;5;220;48;5;101m▓\033[38;5;178;48;5;95m▒\033[38;5;178;48;5;58m▒\033[38;5;178;48;5;95m▒\033[38;5;220;48;5;101m▓\033[38;5;33;48;5;101m▒\033[38;5;50;48;5;137m░\033[38;5;50;48;5;181m▒\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;230m░\033[38;5;117;48;5;144m░\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;180;48;5;58m▒\033[38;5;119;48;5;95m░\033[38;5;50;48;5;247m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▒\033[38;5;131;48;5;236m▒\033[38;5;131;48;5;236m▒\033[38;5;131;48;5;236m▒\033[38;5;131;48;5;236m▒\033[38;5;204;48;5;236m▒\033[38;5;204;48;5;237m▒\033[38;5;204;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;87;48;5;224m░\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;220;48;5;95m▒\033[38;5;50;48;5;247m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;246m▓\033[38;5;50;48;5;181m░\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;172;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;130;48;5;58m░\033[38;5;208;48;5;58m▒\033[38;5;43;48;5;101m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;50;48;5;245m▓\033[38;5;84;48;5;180m░\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m░\033[38;5;130;48;5;94m░\033[38;5;172;48;5;58m░\033[38;5;119;48;5;239m░\033[38;5;50;48;5;144m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m░\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;94;48;5;95m░\033[38;5;209;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▒\033[38;5;80;48;5;187m░\033[38;5;136;48;5;144m▓\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;43;48;5;138m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;187m▒\033[38;5;136;48;5;144m▓\033[38;5;214;48;5;137m▓\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;179m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;94m░\033[38;5;19;48;5;94m░\033[38;5;50;48;5;181m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;174;48;5;236m▒\033[38;5;80;48;5;246m░\033[38;5;179;48;5;101m▓\033[38;5;172;48;5;137m▓\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;101m▒\033[38;5;172;48;5;95m▒\033[38;5;179;48;5;95m▒\033[38;5;214;48;5;95m▒\033[38;5;50;48;5;101m░\033[38;5;1;48;5;16m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;80;48;5;244m▒\033[38;5;214;48;5;238m▓\033[38;5;179;48;5;95m▓\033[38;5;94;48;5;240m▒\033[38;5;94;48;5;95m▓\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;95m▓\033[38;5;34;48;5;237m░\033[38;5;80;48;5;59m░\033[38;5;116;48;5;250m▒\033[38;5;138;48;5;238m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
            $display("\033[0m");

			$display("\nThere is some bug in your code. Errors exceed 100.\n");
			$finish;
		end
	end

endmodule
	
	
		


