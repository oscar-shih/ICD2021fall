`timescale 1ns/1ps

module mode_max(mode, i0, i1, i2, i3, i4);
//DO NOT CHANGE!
	input  [3:0] i0, i1, i2, i3, i4;
	output [3:0] mode;
//---------------------------------------------------
	wire [15:0] a0
	wire [15:0] a1
	wire [15:0] a2
	wire [15:0] a3
	wire [15:0] a4
	
	
endmodule
